`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//
// Montek Singh
// Oct 5, 2021
//
// PLEASE README!
// ==============
//
// This is a self-checking tester for your VGA display driver.
//
// Use this tester carefully!  The names of your top-level input/output
// and internal signals may be different, so some modifications to the tester
// will ne needed.  Here's how to do so:
//
// (1) If the name of an input/output signal in the top-level module is
// different, simply edit the "uut" instantiation block to rename the port name
// to match the name used in the module declaration.  For example, if the "red", "green"
// and "blue" outputs in your top module are instead called "R", "G" and "B",
// change the appropriate line in the "uut" instantiation block:
// FROM
//            .red(red), .green(green), .blue(blue),
// TO
//            .R(red), .G(green), .B(blue),
//
// (2) If the name of an internal signal in the top module is different, simply
// edit the name in the block laeled "INTERNAL SIGNALS".  For example, the tester assumes
// that the vgadisplaydriver instance is called "display", and the x-coordinate within it
// is called "x" (lowercase).  Now suppose your design labels the vgadisplaydriver instance
// as "VGA", and the x-coordinate is labeled uppercase "X".  Then, change the appropriate line
// FROM
//             wire [`xbits-1:0] x = uut.display.x;
// TO
//             wire [`xbits-1:0] x = uut.VGA.X;

// Also, the parameters specifying the names of the
// memory initialization files must match the actual file names.
//
//
// Finally, note that in my bitmap memory, each 12-bit color is encoded as
// RRRRGGGGBBBB (i.e., red is most significant).  If you have chosen a different
// order for the red/green/blue color values, you may see ERROR signals for the
// colors light up.
//
//////////////////////////////////////////////////////////////////////////////////

`include "display640x480.vh"

module tester_sprites_display;

    // Parameters
    localparam Nchars = 64;
    localparam smem_size=1200;              // smem size, 30 rows x 40 cols
    localparam smem_init="screenmem.mem"; 	// text file to initialize screen memory
    localparam bmem_init="bitmapmem.mem"; 	// text file to initialize bitmap memory
    // Parameters derived from above parameters
    localparam charcode_size = $clog2(Nchars);
    localparam bmem_size = Nchars * 256;
     
    // Inputs
    logic clk;

    // Outputs from the top-level display module
    wire hsync, vsync;
    wire [3:0] red, green, blue;
    
    
    // INTERNAL SIGNALS
    // Let's peek inside the top module to check a few signals
    wire [`xbits-1:0] x                    = uut.display.x;
    wire [`ybits-1:0] y                    = uut.display.y;
    wire [$clog2(bmem_size)-1:0] bmem_addr = uut.display.bmem_addr;
    wire [11:0] bmem_color                 = uut.display.bmem_color;
    wire [$clog2(smem_size)-1:0] smem_addr = uut.smem_addr;    // address from vgadisplaydriver to access screen mem
    wire [charcode_size-1:0] charcode      = uut.charcode;     // character code returned by screen mem    
    

    // Instantiate the Unit Under Test (UUT)
    top #(
      .Nchars(Nchars),                    // number of characters/sprites
      .smem_size(smem_size),
      .smem_init(smem_init),
      .bmem_init(bmem_init)
    ) uut(
      .clk(clk), 
      .red(red), .green(green), .blue(blue),
      .hsync(hsync), .vsync(vsync)
    );

//
// CHECK ALL VALUES ABOVE THIS LINE
// YOU SHOULD NOT NEED TO MODIFY ANYTHING BELOW
//

   initial begin
      clk = 0;
      #0.5 clk = 0;
      forever
         #0.5 clk = ~clk;
   end
   
   
   
    // SELF-CHECKING CODE
   
    selfcheck #(.Nchars(Nchars), .smem_size(smem_size)) c();

    wire [$clog2(smem_size)-1:0] c_smem_addr=c.smem_addr;
    wire [$clog2(Nchars)-1:0]  c_charcode=c.charcode;
    wire        c_hsync=c.hsync;
    wire        c_vsync=c.vsync;
    wire [3:0]  c_red=c.red;
    wire [3:0]  c_green=c.green;
    wire [3:0]  c_blue=c.blue;
    wire [`xbits-1:0]  c_x=c.x;
    wire [`ybits-1:0]  c_y=c.y;
    wire [$clog2(Nchars * 256)-1:0] c_bmem_addr=c.bmem_addr;

  
    function mismatch;  // some trickery needed to match two values with don't cares
        input p, q;      // mismatch in a bit position is ignored if q has an 'x' in that bit
        integer p, q;
        mismatch = (((p ^ q) ^ q) !== q);
    endfunction

    wire ERROR;
    wire ERROR_smem_addr      = mismatch(smem_addr, c.smem_addr) ? 1'bx : 1'b0;
    wire ERROR_charcode       = mismatch(charcode, c.charcode) ? 1'bx : 1'b0;
    wire ERROR_hsync          = mismatch(hsync, c.hsync) ? 1'bx : 1'b0;
    wire ERROR_vsync          = mismatch(vsync, c.vsync) ? 1'bx : 1'b0;
    wire ERROR_red            = mismatch(red, c.red) ? 1'bx : 1'b0;
    wire ERROR_green          = mismatch(green, c.green) ? 1'bx : 1'b0;
    wire ERROR_blue           = mismatch(blue, c.blue) ? 1'bx : 1'b0;
    wire ERROR_x              = mismatch(x, c.x) ? 1'bx : 1'b0;
    wire ERROR_y              = mismatch(y, c.y) ? 1'bx : 1'b0;
    wire ERROR_bmem_addr      = mismatch(bmem_addr, c.bmem_addr) ? 1'bx : 1'b0;

    assign ERROR = ERROR_smem_addr | ERROR_charcode | ERROR_hsync | ERROR_vsync
              | ERROR_red | ERROR_green | ERROR_blue
              | ERROR_x | ERROR_y | ERROR_bmem_addr;


    //integer f;
    initial begin
      //f = $fopen("C:/Users/montek/Desktop/output.txt");
      //$fmonitor(f, "#%02d {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h%h, 6'h%h, 1'b%b, 1'b%b, 4'h%h, 4'h%h, 4'h%h, 10'h%h, 10'h%h, 14'h%h};",
      //              $time, smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr);
      #1680000 
      //$fclose(f);
      $finish;
    end

endmodule



// CHECKER MODULE

module selfcheck #(
    parameter Nchars = 4,
    parameter smem_size=1200
)( );
    
    logic [$clog2(smem_size)-1:0] smem_addr;
    logic [$clog2(Nchars)-1:0] charcode;
    logic hsync;
    logic vsync;
    logic [3:0] red;
    logic [3:0] green;
    logic [3:0] blue;
    logic [`xbits-1:0] x;
    logic [`ybits-1:0] y;
    logic [$clog2(Nchars * 256)-1:0] bmem_addr;
    
initial begin
fork


#00 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h000, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h000, 10'h000, 14'h0000};
#04 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#404 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h006, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h065, 10'h000, 14'h0005};
#408 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#808 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h00c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ca, 10'h000, 14'h000a};
#812 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1212 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h012, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h12f, 10'h000, 14'h000f};
#1216 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1616 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h019, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h194, 10'h000, 14'h0004};
#1620 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#2020 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h01f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1f9, 10'h000, 14'h0009};
#2024 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#2424 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h025, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h25e, 10'h000, 14'h000e};
#2428 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#2828 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02c, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2c3, 10'h000, 14'h0003};
#2832 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#3232 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h000, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h008, 10'h001, 14'h0018};
#3236 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#3636 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h006, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h06d, 10'h001, 14'h001d};
#3640 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#4040 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h00d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d2, 10'h001, 14'h0012};
#4044 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#4444 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h013, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h137, 10'h001, 14'h0017};
#4448 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#4848 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h019, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h19c, 10'h001, 14'h001c};
#4852 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#5252 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h020, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h201, 10'h001, 14'h0011};
#5256 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#5656 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h026, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h266, 10'h001, 14'h0016};
#5660 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#6060 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02c, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2cb, 10'h001, 14'h001b};
#6064 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#6464 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h001, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h010, 10'h002, 14'h0020};
#6468 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#6868 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h007, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h075, 10'h002, 14'h0025};
#6872 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#7272 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h00d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0da, 10'h002, 14'h002a};
#7276 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#7676 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h013, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h13f, 10'h002, 14'h002f};
#7680 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#8080 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h01a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1a4, 10'h002, 14'h0024};
#8084 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#8484 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h020, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h209, 10'h002, 14'h0029};
#8488 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#8888 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h026, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h26e, 10'h002, 14'h002e};
#8892 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#9292 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02d, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2d3, 10'h002, 14'h0023};
#9296 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#9696 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h001, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h018, 10'h003, 14'h0038};
#9700 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#10100 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h007, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h07d, 10'h003, 14'h003d};
#10104 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#10504 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h00e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e2, 10'h003, 14'h0032};
#10508 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#10908 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h014, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h147, 10'h003, 14'h0037};
#10912 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#11312 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h01a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1ac, 10'h003, 14'h003c};
#11316 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#11716 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h021, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h211, 10'h003, 14'h0031};
#11720 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#12120 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h027, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h276, 10'h003, 14'h0036};
#12124 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#12524 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02d, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2db, 10'h003, 14'h003b};
#12528 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#12928 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h002, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h020, 10'h004, 14'h0040};
#12932 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#13332 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h008, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h085, 10'h004, 14'h0045};
#13336 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#13736 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h00e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ea, 10'h004, 14'h004a};
#13740 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#14140 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h014, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h14f, 10'h004, 14'h004f};
#14144 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#14544 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h01b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1b4, 10'h004, 14'h0044};
#14548 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#14948 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h021, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h219, 10'h004, 14'h0049};
#14952 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#15352 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h027, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h27e, 10'h004, 14'h004e};
#15356 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#15756 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02e, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2e3, 10'h004, 14'h0043};
#15760 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#16160 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h002, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h028, 10'h005, 14'h0058};
#16164 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#16564 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h008, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h08d, 10'h005, 14'h005d};
#16568 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#16968 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h00f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0f2, 10'h005, 14'h0052};
#16972 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#17372 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h015, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h157, 10'h005, 14'h0057};
#17376 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#17776 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h01b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1bc, 10'h005, 14'h005c};
#17780 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#18180 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h022, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h221, 10'h005, 14'h0051};
#18184 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#18584 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h028, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h286, 10'h005, 14'h0056};
#18588 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#18988 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02e, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2eb, 10'h005, 14'h005b};
#18992 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#19392 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h003, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h030, 10'h006, 14'h0060};
#19396 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#19796 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h009, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h095, 10'h006, 14'h0065};
#19800 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#20200 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h00f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0fa, 10'h006, 14'h006a};
#20204 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#20604 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h015, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h15f, 10'h006, 14'h006f};
#20608 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#21008 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h01c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1c4, 10'h006, 14'h0064};
#21012 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#21412 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h022, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h229, 10'h006, 14'h0069};
#21416 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#21816 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h028, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h28e, 10'h006, 14'h006e};
#21820 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#22220 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02f, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2f3, 10'h006, 14'h0063};
#22224 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#22624 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h003, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h038, 10'h007, 14'h0078};
#22628 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#23028 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h009, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h09d, 10'h007, 14'h007d};
#23032 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#23432 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h010, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h102, 10'h007, 14'h0072};
#23436 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#23836 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h016, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h167, 10'h007, 14'h0077};
#23840 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#24240 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h01c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1cc, 10'h007, 14'h007c};
#24244 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#24644 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h023, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h231, 10'h007, 14'h0071};
#24648 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#25048 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h029, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h296, 10'h007, 14'h0076};
#25052 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#25452 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02f, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2fb, 10'h007, 14'h007b};
#25456 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#25856 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h004, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h040, 10'h008, 14'h0080};
#25860 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#26260 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h00a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0a5, 10'h008, 14'h0085};
#26264 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#26664 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h010, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h10a, 10'h008, 14'h008a};
#26668 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#27068 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h016, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h16f, 10'h008, 14'h008f};
#27072 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#27472 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h01d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1d4, 10'h008, 14'h0084};
#27476 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#27876 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h023, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h239, 10'h008, 14'h0089};
#27880 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#28280 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h029, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h29e, 10'h008, 14'h008e};
#28284 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#28684 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h030, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h303, 10'h008, 14'h0083};
#28688 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#29088 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h004, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h048, 10'h009, 14'h0098};
#29092 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#29492 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h00a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ad, 10'h009, 14'h009d};
#29496 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#29896 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h011, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h112, 10'h009, 14'h0092};
#29900 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#30300 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h017, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h177, 10'h009, 14'h0097};
#30304 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#30704 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h01d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1dc, 10'h009, 14'h009c};
#30708 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#31108 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h024, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h241, 10'h009, 14'h0091};
#31112 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#31512 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02a, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2a6, 10'h009, 14'h0096};
#31516 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#31916 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h030, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h30b, 10'h009, 14'h009b};
#31920 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#32320 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h005, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h050, 10'h00a, 14'h00a0};
#32324 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#32724 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h00b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0b5, 10'h00a, 14'h00a5};
#32728 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#33128 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h011, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h11a, 10'h00a, 14'h00aa};
#33132 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#33532 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h017, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h17f, 10'h00a, 14'h00af};
#33536 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#33936 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h01e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1e4, 10'h00a, 14'h00a4};
#33940 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#34340 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h024, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h249, 10'h00a, 14'h00a9};
#34344 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#34744 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02a, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2ae, 10'h00a, 14'h00ae};
#34748 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#35148 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h031, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h313, 10'h00a, 14'h00a3};
#35152 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#35552 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h005, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h058, 10'h00b, 14'h00b8};
#35556 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#35956 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h00b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0bd, 10'h00b, 14'h00bd};
#35960 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#36360 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h012, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h122, 10'h00b, 14'h00b2};
#36364 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#36764 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h018, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h187, 10'h00b, 14'h00b7};
#36768 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#37168 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h01e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1ec, 10'h00b, 14'h00bc};
#37172 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#37572 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h025, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h251, 10'h00b, 14'h00b1};
#37576 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#37976 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02b, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2b6, 10'h00b, 14'h00b6};
#37980 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#38380 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h031, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h31b, 10'h00b, 14'h00bb};
#38384 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#38784 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h006, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h060, 10'h00c, 14'h00c0};
#38788 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#39188 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h00c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c5, 10'h00c, 14'h00c5};
#39192 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#39592 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h012, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h12a, 10'h00c, 14'h00ca};
#39596 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#39996 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h018, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h18f, 10'h00c, 14'h00cf};
#40000 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#40400 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h01f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1f4, 10'h00c, 14'h00c4};
#40404 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#40804 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h025, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h259, 10'h00c, 14'h00c9};
#40808 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#41208 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02b, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2be, 10'h00c, 14'h00ce};
#41212 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#41612 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h000, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h003, 10'h00d, 14'h00d3};
#41616 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#42016 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h006, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h068, 10'h00d, 14'h00d8};
#42020 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#42420 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h00c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0cd, 10'h00d, 14'h00dd};
#42424 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#42824 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h013, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h132, 10'h00d, 14'h00d2};
#42828 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#43228 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h019, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h197, 10'h00d, 14'h00d7};
#43232 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#43632 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h01f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1fc, 10'h00d, 14'h00dc};
#43636 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#44036 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h026, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h261, 10'h00d, 14'h00d1};
#44040 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#44440 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02c, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2c6, 10'h00d, 14'h00d6};
#44444 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#44844 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h000, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00b, 10'h00e, 14'h00eb};
#44848 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#45248 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h007, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h070, 10'h00e, 14'h00e0};
#45252 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#45652 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h00d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d5, 10'h00e, 14'h00e5};
#45656 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#46056 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h013, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h13a, 10'h00e, 14'h00ea};
#46060 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#46460 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h019, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h19f, 10'h00e, 14'h00ef};
#46464 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#46864 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h020, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h204, 10'h00e, 14'h00e4};
#46868 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#47268 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h026, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h269, 10'h00e, 14'h00e9};
#47272 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#47672 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02c, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2ce, 10'h00e, 14'h00ee};
#47676 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#48076 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h001, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h013, 10'h00f, 14'h00f3};
#48080 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#48480 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h007, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h078, 10'h00f, 14'h00f8};
#48484 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#48884 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h00d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0dd, 10'h00f, 14'h00fd};
#48888 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#49288 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h014, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h142, 10'h00f, 14'h00f2};
#49292 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#49692 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h01a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1a7, 10'h00f, 14'h00f7};
#49696 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#50096 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h020, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h20c, 10'h00f, 14'h00fc};
#50100 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#50500 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h027, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h271, 10'h00f, 14'h00f1};
#50504 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#50904 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02d, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2d6, 10'h00f, 14'h00f6};
#50908 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#51308 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h029, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h01b, 10'h010, 14'h000b};
#51312 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#51712 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h030, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h080, 10'h010, 14'h0000};
#51716 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#52116 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h036, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e5, 10'h010, 14'h0005};
#52120 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#52520 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h03c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h14a, 10'h010, 14'h000a};
#52524 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#52924 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h042, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1af, 10'h010, 14'h000f};
#52928 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#53328 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h049, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h214, 10'h010, 14'h0004};
#53332 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#53732 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h04f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h279, 10'h010, 14'h0009};
#53736 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#54136 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h055, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2de, 10'h010, 14'h000e};
#54140 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#54540 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h023, 10'h011, 14'h0013};
#54544 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#54944 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h030, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h088, 10'h011, 14'h0018};
#54948 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#55348 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h036, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ed, 10'h011, 14'h001d};
#55352 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#55752 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h03d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h152, 10'h011, 14'h0012};
#55756 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#56156 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h043, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1b7, 10'h011, 14'h0017};
#56160 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#56560 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h049, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h21c, 10'h011, 14'h001c};
#56564 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#56964 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h050, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h281, 10'h011, 14'h0011};
#56968 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#57368 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h056, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2e6, 10'h011, 14'h0016};
#57372 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#57772 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02b, 10'h012, 14'h002b};
#57776 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#58176 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h031, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h090, 10'h012, 14'h0020};
#58180 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#58580 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h037, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0f5, 10'h012, 14'h0025};
#58584 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#58984 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h03d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h15a, 10'h012, 14'h002a};
#58988 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#59388 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h043, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1bf, 10'h012, 14'h002f};
#59392 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#59792 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h04a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h224, 10'h012, 14'h0024};
#59796 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#60196 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h050, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h289, 10'h012, 14'h0029};
#60200 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#60600 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h056, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2ee, 10'h012, 14'h002e};
#60604 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#61004 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h033, 10'h013, 14'h0033};
#61008 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#61408 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h031, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h098, 10'h013, 14'h0038};
#61412 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#61812 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h037, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0fd, 10'h013, 14'h003d};
#61816 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#62216 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h03e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h162, 10'h013, 14'h0032};
#62220 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#62620 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h044, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1c7, 10'h013, 14'h0037};
#62624 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#63024 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h04a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h22c, 10'h013, 14'h003c};
#63028 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#63428 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h051, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h291, 10'h013, 14'h0031};
#63432 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#63832 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h057, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2f6, 10'h013, 14'h0036};
#63836 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#64236 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h03b, 10'h014, 14'h004b};
#64240 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#64640 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h032, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0a0, 10'h014, 14'h0040};
#64644 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#65044 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h038, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h105, 10'h014, 14'h0045};
#65048 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#65448 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h03e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h16a, 10'h014, 14'h004a};
#65452 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#65852 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h044, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1cf, 10'h014, 14'h004f};
#65856 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#66256 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h04b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h234, 10'h014, 14'h0044};
#66260 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#66660 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h051, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h299, 10'h014, 14'h0049};
#66664 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#67064 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h057, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2fe, 10'h014, 14'h004e};
#67068 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#67468 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h043, 10'h015, 14'h0053};
#67472 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#67872 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h032, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0a8, 10'h015, 14'h0058};
#67876 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#68276 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h038, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h10d, 10'h015, 14'h005d};
#68280 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#68680 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h03f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h172, 10'h015, 14'h0052};
#68684 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#69084 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h045, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1d7, 10'h015, 14'h0057};
#69088 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#69488 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h04b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h23c, 10'h015, 14'h005c};
#69492 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#69892 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h052, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2a1, 10'h015, 14'h0051};
#69896 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#70296 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h058, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h306, 10'h015, 14'h0056};
#70300 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#70700 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h04b, 10'h016, 14'h006b};
#70704 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#71104 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h033, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0b0, 10'h016, 14'h0060};
#71108 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#71508 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h039, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h115, 10'h016, 14'h0065};
#71512 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#71912 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h03f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h17a, 10'h016, 14'h006a};
#71916 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#72316 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h045, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1df, 10'h016, 14'h006f};
#72320 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#72720 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h04c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h244, 10'h016, 14'h0064};
#72724 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#73124 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h052, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2a9, 10'h016, 14'h0069};
#73128 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#73528 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h058, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h30e, 10'h016, 14'h006e};
#73532 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#73932 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h053, 10'h017, 14'h0073};
#73936 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#74336 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h033, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0b8, 10'h017, 14'h0078};
#74340 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#74740 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h039, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h11d, 10'h017, 14'h007d};
#74744 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#75144 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h040, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h182, 10'h017, 14'h0072};
#75148 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#75548 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h046, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1e7, 10'h017, 14'h0077};
#75552 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#75952 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h04c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h24c, 10'h017, 14'h007c};
#75956 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#76356 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h053, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2b1, 10'h017, 14'h0071};
#76360 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#76760 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h059, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h316, 10'h017, 14'h0076};
#76764 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#77164 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h05b, 10'h018, 14'h008b};
#77168 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#77568 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h034, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c0, 10'h018, 14'h0080};
#77572 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#77972 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h03a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h125, 10'h018, 14'h0085};
#77976 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#78376 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h040, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h18a, 10'h018, 14'h008a};
#78380 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#78780 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h046, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1ef, 10'h018, 14'h008f};
#78784 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#79184 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h04d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h254, 10'h018, 14'h0084};
#79188 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#79588 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h053, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2b9, 10'h018, 14'h0089};
#79592 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#79992 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h059, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h31e, 10'h018, 14'h008e};
#79996 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#80396 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h063, 10'h019, 14'h0093};
#80400 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#80800 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h034, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c8, 10'h019, 14'h0098};
#80804 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#81204 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h03a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h12d, 10'h019, 14'h009d};
#81208 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#81608 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h041, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h192, 10'h019, 14'h0092};
#81612 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#82012 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h047, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1f7, 10'h019, 14'h0097};
#82016 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#82416 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h04d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h25c, 10'h019, 14'h009c};
#82420 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#82820 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h054, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2c1, 10'h019, 14'h0091};
#82824 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#83224 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h028, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h006, 10'h01a, 14'h00a6};
#83228 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#83628 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h06b, 10'h01a, 14'h00ab};
#83632 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#84032 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h035, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d0, 10'h01a, 14'h00a0};
#84036 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#84436 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h03b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h135, 10'h01a, 14'h00a5};
#84440 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#84840 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h041, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h19a, 10'h01a, 14'h00aa};
#84844 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#85244 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h047, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1ff, 10'h01a, 14'h00af};
#85248 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#85648 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h04e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h264, 10'h01a, 14'h00a4};
#85652 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#86052 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h054, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2c9, 10'h01a, 14'h00a9};
#86056 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#86456 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h028, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00e, 10'h01b, 14'h00be};
#86460 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#86860 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h073, 10'h01b, 14'h00b3};
#86864 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#87264 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h035, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d8, 10'h01b, 14'h00b8};
#87268 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#87668 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h03b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h13d, 10'h01b, 14'h00bd};
#87672 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#88072 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h042, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1a2, 10'h01b, 14'h00b2};
#88076 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#88476 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h048, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h207, 10'h01b, 14'h00b7};
#88480 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#88880 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h04e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h26c, 10'h01b, 14'h00bc};
#88884 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#89284 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h055, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2d1, 10'h01b, 14'h00b1};
#89288 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#89688 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h029, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h016, 10'h01c, 14'h00c6};
#89692 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#90092 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h07b, 10'h01c, 14'h00cb};
#90096 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#90496 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h036, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e0, 10'h01c, 14'h00c0};
#90500 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#90900 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h03c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h145, 10'h01c, 14'h00c5};
#90904 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#91304 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h042, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1aa, 10'h01c, 14'h00ca};
#91308 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#91708 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h048, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h20f, 10'h01c, 14'h00cf};
#91712 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#92112 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h04f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h274, 10'h01c, 14'h00c4};
#92116 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#92516 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h055, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2d9, 10'h01c, 14'h00c9};
#92520 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#92920 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h029, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h01e, 10'h01d, 14'h00de};
#92924 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#93324 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h030, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h083, 10'h01d, 14'h00d3};
#93328 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#93728 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h036, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e8, 10'h01d, 14'h00d8};
#93732 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#94132 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h03c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h14d, 10'h01d, 14'h00dd};
#94136 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#94536 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h043, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1b2, 10'h01d, 14'h00d2};
#94540 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#94940 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h049, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h217, 10'h01d, 14'h00d7};
#94944 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#95344 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h04f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h27c, 10'h01d, 14'h00dc};
#95348 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#95748 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h056, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2e1, 10'h01d, 14'h00d1};
#95752 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#96152 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h026, 10'h01e, 14'h00e6};
#96156 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#96556 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h030, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h08b, 10'h01e, 14'h00eb};
#96560 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#96960 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h037, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0f0, 10'h01e, 14'h00e0};
#96964 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#97364 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h03d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h155, 10'h01e, 14'h00e5};
#97368 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#97768 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h043, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1ba, 10'h01e, 14'h00ea};
#97772 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#98172 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h049, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h21f, 10'h01e, 14'h00ef};
#98176 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#98576 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h050, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h284, 10'h01e, 14'h00e4};
#98580 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#98980 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h056, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2e9, 10'h01e, 14'h00e9};
#98984 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#99384 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h02a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02e, 10'h01f, 14'h00fe};
#99388 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#99788 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h031, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h093, 10'h01f, 14'h00f3};
#99792 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#100192 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h037, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0f8, 10'h01f, 14'h00f8};
#100196 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#100596 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h03d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h15d, 10'h01f, 14'h00fd};
#100600 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#101000 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h044, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1c2, 10'h01f, 14'h00f2};
#101004 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#101404 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h04a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h227, 10'h01f, 14'h00f7};
#101408 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#101808 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h050, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h28c, 10'h01f, 14'h00fc};
#101812 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#102212 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h057, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2f1, 10'h01f, 14'h00f1};
#102216 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#102616 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h053, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h036, 10'h020, 14'h0006};
#102620 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#103020 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h059, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h09b, 10'h020, 14'h000b};
#103024 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#103424 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h060, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h100, 10'h020, 14'h0000};
#103428 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#103828 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h066, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h165, 10'h020, 14'h0005};
#103832 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#104232 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h06c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1ca, 10'h020, 14'h000a};
#104236 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#104636 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h072, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h22f, 10'h020, 14'h000f};
#104640 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#105040 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h079, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h294, 10'h020, 14'h0004};
#105044 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#105444 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07f, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2f9, 10'h020, 14'h0009};
#105448 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#105848 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h053, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h03e, 10'h021, 14'h001e};
#105852 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#106252 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h05a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0a3, 10'h021, 14'h0013};
#106256 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#106656 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h060, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h108, 10'h021, 14'h0018};
#106660 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#107060 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h066, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h16d, 10'h021, 14'h001d};
#107064 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#107464 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h06d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1d2, 10'h021, 14'h0012};
#107468 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#107868 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h073, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h237, 10'h021, 14'h0017};
#107872 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#108272 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h079, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h29c, 10'h021, 14'h001c};
#108276 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#108676 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h080, 6'h01, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h301, 10'h021, 14'h0111};
#108680 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#109080 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h054, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h046, 10'h022, 14'h0026};
#109084 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#109484 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h05a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ab, 10'h022, 14'h002b};
#109488 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#109888 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h061, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h110, 10'h022, 14'h0020};
#109892 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#110292 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h067, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h175, 10'h022, 14'h0025};
#110296 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#110696 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h06d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1da, 10'h022, 14'h002a};
#110700 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#111100 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h073, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h23f, 10'h022, 14'h002f};
#111104 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#111504 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07a, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2a4, 10'h022, 14'h0024};
#111508 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#111908 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h080, 6'h01, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h309, 10'h022, 14'h0129};
#111912 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#112312 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h054, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h04e, 10'h023, 14'h003e};
#112316 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#112716 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h05b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0b3, 10'h023, 14'h0033};
#112720 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#113120 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h061, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h118, 10'h023, 14'h0038};
#113124 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#113524 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h067, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h17d, 10'h023, 14'h003d};
#113528 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#113928 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h06e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1e2, 10'h023, 14'h0032};
#113932 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#114332 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h074, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h247, 10'h023, 14'h0037};
#114336 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#114736 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07a, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2ac, 10'h023, 14'h003c};
#114740 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#115140 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h081, 6'h01, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h311, 10'h023, 14'h0131};
#115144 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#115544 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h055, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h056, 10'h024, 14'h0046};
#115548 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#115948 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h05b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0bb, 10'h024, 14'h004b};
#115952 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#116352 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h062, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h120, 10'h024, 14'h0040};
#116356 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#116756 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h068, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h185, 10'h024, 14'h0045};
#116760 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#117160 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h06e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1ea, 10'h024, 14'h004a};
#117164 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#117564 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h074, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h24f, 10'h024, 14'h004f};
#117568 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#117968 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07b, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2b4, 10'h024, 14'h0044};
#117972 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#118372 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h081, 6'h01, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h319, 10'h024, 14'h0149};
#118376 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#118776 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h055, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h05e, 10'h025, 14'h005e};
#118780 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#119180 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h05c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c3, 10'h025, 14'h0053};
#119184 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#119584 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h062, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h128, 10'h025, 14'h0058};
#119588 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#119988 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h068, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h18d, 10'h025, 14'h005d};
#119992 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#120392 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h06f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1f2, 10'h025, 14'h0052};
#120396 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#120796 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h075, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h257, 10'h025, 14'h0057};
#120800 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#121200 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07b, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2bc, 10'h025, 14'h005c};
#121204 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#121604 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h050, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h001, 10'h026, 14'h0061};
#121608 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#122008 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h056, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h066, 10'h026, 14'h0066};
#122012 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#122412 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h05c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0cb, 10'h026, 14'h006b};
#122416 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#122816 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h063, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h130, 10'h026, 14'h0060};
#122820 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#123220 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h069, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h195, 10'h026, 14'h0065};
#123224 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#123624 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h06f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1fa, 10'h026, 14'h006a};
#123628 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#124028 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h075, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h25f, 10'h026, 14'h006f};
#124032 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#124432 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07c, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2c4, 10'h026, 14'h0064};
#124436 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#124836 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h050, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h009, 10'h027, 14'h0079};
#124840 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#125240 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h056, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h06e, 10'h027, 14'h007e};
#125244 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#125644 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h05d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d3, 10'h027, 14'h0073};
#125648 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#126048 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h063, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h138, 10'h027, 14'h0078};
#126052 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#126452 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h069, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h19d, 10'h027, 14'h007d};
#126456 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#126856 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h070, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h202, 10'h027, 14'h0072};
#126860 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#127260 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h076, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h267, 10'h027, 14'h0077};
#127264 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#127664 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07c, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2cc, 10'h027, 14'h007c};
#127668 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#128068 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h051, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h011, 10'h028, 14'h0081};
#128072 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#128472 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h057, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h076, 10'h028, 14'h0086};
#128476 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#128876 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h05d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0db, 10'h028, 14'h008b};
#128880 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#129280 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h064, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h140, 10'h028, 14'h0080};
#129284 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#129684 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h06a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1a5, 10'h028, 14'h0085};
#129688 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#130088 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h070, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h20a, 10'h028, 14'h008a};
#130092 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#130492 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h076, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h26f, 10'h028, 14'h008f};
#130496 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#130896 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07d, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2d4, 10'h028, 14'h0084};
#130900 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#131300 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h051, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h019, 10'h029, 14'h0099};
#131304 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#131704 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h057, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h07e, 10'h029, 14'h009e};
#131708 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#132108 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h05e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e3, 10'h029, 14'h0093};
#132112 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#132512 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h064, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h148, 10'h029, 14'h0098};
#132516 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#132916 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h06a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1ad, 10'h029, 14'h009d};
#132920 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#133320 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h071, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h212, 10'h029, 14'h0092};
#133324 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#133724 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h077, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h277, 10'h029, 14'h0097};
#133728 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#134128 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07d, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2dc, 10'h029, 14'h009c};
#134132 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#134532 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h052, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h021, 10'h02a, 14'h00a1};
#134536 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#134936 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h058, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h086, 10'h02a, 14'h00a6};
#134940 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#135340 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h05e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0eb, 10'h02a, 14'h00ab};
#135344 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#135744 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h065, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h150, 10'h02a, 14'h00a0};
#135748 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#136148 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h06b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1b5, 10'h02a, 14'h00a5};
#136152 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#136552 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h071, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h21a, 10'h02a, 14'h00aa};
#136556 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#136956 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h077, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h27f, 10'h02a, 14'h00af};
#136960 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#137360 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07e, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2e4, 10'h02a, 14'h00a4};
#137364 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#137764 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h052, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h029, 10'h02b, 14'h00b9};
#137768 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#138168 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h058, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h08e, 10'h02b, 14'h00be};
#138172 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#138572 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h05f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0f3, 10'h02b, 14'h00b3};
#138576 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#138976 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h065, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h158, 10'h02b, 14'h00b8};
#138980 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#139380 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h06b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1bd, 10'h02b, 14'h00bd};
#139384 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#139784 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h072, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h222, 10'h02b, 14'h00b2};
#139788 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#140188 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h078, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h287, 10'h02b, 14'h00b7};
#140192 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#140592 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07e, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2ec, 10'h02b, 14'h00bc};
#140596 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#140996 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h053, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h031, 10'h02c, 14'h00c1};
#141000 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#141400 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h059, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h096, 10'h02c, 14'h00c6};
#141404 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#141804 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h05f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0fb, 10'h02c, 14'h00cb};
#141808 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#142208 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h066, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h160, 10'h02c, 14'h00c0};
#142212 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#142612 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h06c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1c5, 10'h02c, 14'h00c5};
#142616 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#143016 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h072, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h22a, 10'h02c, 14'h00ca};
#143020 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#143420 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h078, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h28f, 10'h02c, 14'h00cf};
#143424 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#143824 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07f, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2f4, 10'h02c, 14'h00c4};
#143828 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#144228 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h053, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h039, 10'h02d, 14'h00d9};
#144232 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#144632 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h059, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h09e, 10'h02d, 14'h00de};
#144636 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#145036 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h060, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h103, 10'h02d, 14'h00d3};
#145040 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#145440 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h066, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h168, 10'h02d, 14'h00d8};
#145444 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#145844 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h06c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1cd, 10'h02d, 14'h00dd};
#145848 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#146248 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h073, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h232, 10'h02d, 14'h00d2};
#146252 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#146652 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h079, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h297, 10'h02d, 14'h00d7};
#146656 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#147056 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07f, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2fc, 10'h02d, 14'h00dc};
#147060 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#147460 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h054, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h041, 10'h02e, 14'h00e1};
#147464 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#147864 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h05a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0a6, 10'h02e, 14'h00e6};
#147868 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#148268 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h060, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h10b, 10'h02e, 14'h00eb};
#148272 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#148672 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h067, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h170, 10'h02e, 14'h00e0};
#148676 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#149076 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h06d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1d5, 10'h02e, 14'h00e5};
#149080 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#149480 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h073, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h23a, 10'h02e, 14'h00ea};
#149484 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#149884 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h079, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h29f, 10'h02e, 14'h00ef};
#149888 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#150288 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h080, 6'h01, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h304, 10'h02e, 14'h01e4};
#150292 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#150692 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h054, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h049, 10'h02f, 14'h00f9};
#150696 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#151096 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h05a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ae, 10'h02f, 14'h00fe};
#151100 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#151500 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h061, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h113, 10'h02f, 14'h00f3};
#151504 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#151904 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h067, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h178, 10'h02f, 14'h00f8};
#151908 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#152308 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h06d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1dd, 10'h02f, 14'h00fd};
#152312 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#152712 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h074, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h242, 10'h02f, 14'h00f2};
#152716 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#153116 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07a, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2a7, 10'h02f, 14'h00f7};
#153120 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#153520 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h080, 6'h01, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h30c, 10'h02f, 14'h01fc};
#153524 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#153924 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h051, 10'h030, 14'h0001};
#153928 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#154328 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h083, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0b6, 10'h030, 14'h0006};
#154332 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#154732 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h089, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h11b, 10'h030, 14'h020b};
#154736 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#155136 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h090, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h180, 10'h030, 14'h0000};
#155140 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#155540 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h096, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1e5, 10'h030, 14'h0005};
#155544 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#155944 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h09c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h24a, 10'h030, 14'h000a};
#155948 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#156348 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a2, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2af, 10'h030, 14'h000f};
#156352 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#156752 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a9, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h314, 10'h030, 14'h0004};
#156756 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#157156 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h059, 10'h031, 14'h0019};
#157160 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#157560 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h083, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0be, 10'h031, 14'h001e};
#157564 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#157964 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h08a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h123, 10'h031, 14'h0013};
#157968 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#158368 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h090, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h188, 10'h031, 14'h0018};
#158372 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#158772 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h096, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1ed, 10'h031, 14'h001d};
#158776 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#159176 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h09d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h252, 10'h031, 14'h0012};
#159180 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#159580 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a3, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2b7, 10'h031, 14'h0017};
#159584 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#159984 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a9, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h31c, 10'h031, 14'h001c};
#159988 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#160388 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h061, 10'h032, 14'h0021};
#160392 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#160792 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h084, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c6, 10'h032, 14'h0026};
#160796 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#161196 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h08a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h12b, 10'h032, 14'h002b};
#161200 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#161600 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h091, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h190, 10'h032, 14'h0020};
#161604 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#162004 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h097, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h1f5, 10'h032, 14'h0125};
#162008 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#162408 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h09d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h25a, 10'h032, 14'h002a};
#162412 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#162812 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a3, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2bf, 10'h032, 14'h002f};
#162816 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#163216 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h078, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h004, 10'h033, 14'h0034};
#163220 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#163620 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h069, 10'h033, 14'h0039};
#163624 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#164024 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h084, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ce, 10'h033, 14'h003e};
#164028 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#164428 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h08b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h133, 10'h033, 14'h0033};
#164432 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#164832 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h091, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h198, 10'h033, 14'h0038};
#164836 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#165236 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h097, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h1fd, 10'h033, 14'h013d};
#165240 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#165640 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h09e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h262, 10'h033, 14'h0032};
#165644 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#166044 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a4, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2c7, 10'h033, 14'h0037};
#166048 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#166448 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h078, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00c, 10'h034, 14'h004c};
#166452 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#166852 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h071, 10'h034, 14'h0041};
#166856 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#167256 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h085, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d6, 10'h034, 14'h0046};
#167260 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#167660 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h08b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h13b, 10'h034, 14'h004b};
#167664 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#168064 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h092, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1a0, 10'h034, 14'h0040};
#168068 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#168468 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h098, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h205, 10'h034, 14'h0145};
#168472 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#168872 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h09e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h26a, 10'h034, 14'h004a};
#168876 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#169276 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a4, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2cf, 10'h034, 14'h004f};
#169280 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#169680 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h079, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h014, 10'h035, 14'h0054};
#169684 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#170084 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h079, 10'h035, 14'h0059};
#170088 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#170488 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h085, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0de, 10'h035, 14'h005e};
#170492 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#170892 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h08c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h143, 10'h035, 14'h0053};
#170896 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#171296 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h092, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1a8, 10'h035, 14'h0058};
#171300 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#171700 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h098, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h20d, 10'h035, 14'h015d};
#171704 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#172104 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h09f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h272, 10'h035, 14'h0052};
#172108 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#172508 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a5, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2d7, 10'h035, 14'h0057};
#172512 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#172912 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h079, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h01c, 10'h036, 14'h006c};
#172916 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#173316 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h080, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h081, 10'h036, 14'h0161};
#173320 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#173720 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h086, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e6, 10'h036, 14'h0066};
#173724 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#174124 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h08c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h14b, 10'h036, 14'h006b};
#174128 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#174528 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h093, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1b0, 10'h036, 14'h0060};
#174532 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#174932 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h099, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h215, 10'h036, 14'h0165};
#174936 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#175336 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h09f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h27a, 10'h036, 14'h006a};
#175340 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#175740 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a5, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2df, 10'h036, 14'h006f};
#175744 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#176144 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h024, 10'h037, 14'h0074};
#176148 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#176548 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h080, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h089, 10'h037, 14'h0179};
#176552 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#176952 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h086, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ee, 10'h037, 14'h007e};
#176956 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#177356 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h08d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h153, 10'h037, 14'h0073};
#177360 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#177760 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h093, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1b8, 10'h037, 14'h0078};
#177764 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#178164 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h099, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h21d, 10'h037, 14'h017d};
#178168 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#178568 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a0, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h282, 10'h037, 14'h0072};
#178572 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#178972 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a6, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2e7, 10'h037, 14'h0077};
#178976 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#179376 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02c, 10'h038, 14'h008c};
#179380 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#179780 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h081, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h091, 10'h038, 14'h0181};
#179784 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#180184 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h087, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h0f6, 10'h038, 14'h0286};
#180188 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#180588 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h08d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h15b, 10'h038, 14'h008b};
#180592 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#180992 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h094, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h1c0, 10'h038, 14'h0380};
#180996 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#181396 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h09a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h225, 10'h038, 14'h0085};
#181400 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#181800 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a0, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h28a, 10'h038, 14'h008a};
#181804 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#182204 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a6, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2ef, 10'h038, 14'h008f};
#182208 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#182608 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h034, 10'h039, 14'h0094};
#182612 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#183012 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h081, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h099, 10'h039, 14'h0199};
#183016 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#183416 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h087, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h0fe, 10'h039, 14'h029e};
#183420 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#183820 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h08e, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h163, 10'h039, 14'h0393};
#183824 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#184224 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h094, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h1c8, 10'h039, 14'h0398};
#184228 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#184628 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h09a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h22d, 10'h039, 14'h009d};
#184632 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#185032 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a1, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h292, 10'h039, 14'h0092};
#185036 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#185436 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a7, 6'h01, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2f7, 10'h039, 14'h0197};
#185440 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#185840 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h03c, 10'h03a, 14'h00ac};
#185844 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#186244 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h082, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0a1, 10'h03a, 14'h01a1};
#186248 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#186648 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h088, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h106, 10'h03a, 14'h02a6};
#186652 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#187052 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h08e, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h16b, 10'h03a, 14'h03ab};
#187056 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#187456 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h095, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1d0, 10'h03a, 14'h00a0};
#187460 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#187860 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h09b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h235, 10'h03a, 14'h00a5};
#187864 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#188264 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a1, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h29a, 10'h03a, 14'h00aa};
#188268 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#188668 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a7, 6'h01, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2ff, 10'h03a, 14'h01af};
#188672 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#189072 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h044, 10'h03b, 14'h00b4};
#189076 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#189476 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h082, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0a9, 10'h03b, 14'h01b9};
#189480 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#189880 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h088, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h10e, 10'h03b, 14'h02be};
#189884 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#190284 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h08f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h173, 10'h03b, 14'h00b3};
#190288 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#190688 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h095, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1d8, 10'h03b, 14'h00b8};
#190692 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#191092 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h09b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h23d, 10'h03b, 14'h00bd};
#191096 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#191496 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a2, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2a2, 10'h03b, 14'h00b2};
#191500 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#191900 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a8, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h307, 10'h03b, 14'h00b7};
#191904 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#192304 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h04c, 10'h03c, 14'h00cc};
#192308 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#192708 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h083, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0b1, 10'h03c, 14'h00c1};
#192712 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#193112 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h089, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h116, 10'h03c, 14'h02c6};
#193116 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#193516 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h08f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h17b, 10'h03c, 14'h00cb};
#193520 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#193920 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h096, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1e0, 10'h03c, 14'h00c0};
#193924 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#194324 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h09c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h245, 10'h03c, 14'h00c5};
#194328 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#194728 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a2, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2aa, 10'h03c, 14'h00ca};
#194732 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#195132 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a8, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h30f, 10'h03c, 14'h00cf};
#195136 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#195536 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h054, 10'h03d, 14'h00d4};
#195540 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#195940 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h083, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0b9, 10'h03d, 14'h00d9};
#195944 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#196344 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h089, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h11e, 10'h03d, 14'h02de};
#196348 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#196748 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h090, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h183, 10'h03d, 14'h00d3};
#196752 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#197152 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h096, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1e8, 10'h03d, 14'h00d8};
#197156 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#197556 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h09c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h24d, 10'h03d, 14'h00dd};
#197560 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#197960 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a3, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2b2, 10'h03d, 14'h00d2};
#197964 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#198364 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a9, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h317, 10'h03d, 14'h00d7};
#198368 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#198768 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h05c, 10'h03e, 14'h00ec};
#198772 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#199172 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h084, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c1, 10'h03e, 14'h00e1};
#199176 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#199576 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h08a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h126, 10'h03e, 14'h00e6};
#199580 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#199980 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h090, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h18b, 10'h03e, 14'h00eb};
#199984 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#200384 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h097, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h1f0, 10'h03e, 14'h01e0};
#200388 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#200788 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h09d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h255, 10'h03e, 14'h00e5};
#200792 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#201192 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a3, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2ba, 10'h03e, 14'h00ea};
#201196 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#201596 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a9, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h31f, 10'h03e, 14'h00ef};
#201600 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#202000 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h07e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h064, 10'h03f, 14'h00f4};
#202004 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#202404 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h084, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c9, 10'h03f, 14'h00f9};
#202408 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#202808 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h08a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h12e, 10'h03f, 14'h00fe};
#202812 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#203212 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h091, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h193, 10'h03f, 14'h00f3};
#203216 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#203616 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h097, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h1f8, 10'h03f, 14'h01f8};
#203620 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#204020 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h09d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h25d, 10'h03f, 14'h00fd};
#204024 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#204424 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a4, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2c2, 10'h03f, 14'h00f2};
#204428 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#204828 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h007, 10'h040, 14'h0007};
#204832 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#205232 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a6, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h06c, 10'h040, 14'h000c};
#205236 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#205636 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ad, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d1, 10'h040, 14'h0001};
#205640 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#206040 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0b3, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h136, 10'h040, 14'h0006};
#206044 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#206444 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0b9, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h19b, 10'h040, 14'h000b};
#206448 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#206848 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h200, 10'h040, 14'h0000};
#206852 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#207252 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c6, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h265, 10'h040, 14'h0005};
#207256 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#207656 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0cc, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2ca, 10'h040, 14'h000a};
#207660 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#208060 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00f, 10'h041, 14'h001f};
#208064 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#208464 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a7, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h074, 10'h041, 14'h0114};
#208468 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#208868 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ad, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d9, 10'h041, 14'h0019};
#208872 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#209272 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0b3, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h13e, 10'h041, 14'h001e};
#209276 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#209676 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ba, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1a3, 10'h041, 14'h0013};
#209680 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#210080 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h208, 10'h041, 14'h0018};
#210084 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#210484 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c6, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h26d, 10'h041, 14'h001d};
#210488 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#210888 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0cd, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2d2, 10'h041, 14'h0012};
#210892 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#211292 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h017, 10'h042, 14'h0027};
#211296 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#211696 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a7, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h07c, 10'h042, 14'h012c};
#211700 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#212100 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ae, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h0e1, 10'h042, 14'h0221};
#212104 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#212504 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0b4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h146, 10'h042, 14'h0026};
#212508 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#212908 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ba, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1ab, 10'h042, 14'h002b};
#212912 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#213312 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h210, 10'h042, 14'h0020};
#213316 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#213716 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c7, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h275, 10'h042, 14'h0025};
#213720 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#214120 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0cd, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2da, 10'h042, 14'h002a};
#214124 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#214524 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h01f, 10'h043, 14'h003f};
#214528 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#214928 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a8, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h084, 10'h043, 14'h0034};
#214932 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#215332 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ae, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h0e9, 10'h043, 14'h0239};
#215336 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#215736 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0b4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h14e, 10'h043, 14'h003e};
#215740 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#216140 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0bb, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h1b3, 10'h043, 14'h0333};
#216144 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#216544 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h218, 10'h043, 14'h0038};
#216548 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#216948 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c7, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h27d, 10'h043, 14'h003d};
#216952 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#217352 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ce, 6'h01, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2e2, 10'h043, 14'h0132};
#217356 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#217756 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a2, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h027, 10'h044, 14'h0047};
#217760 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#218160 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a8, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h08c, 10'h044, 14'h004c};
#218164 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#218564 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0af, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0f1, 10'h044, 14'h0041};
#218568 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#218968 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0b5, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h156, 10'h044, 14'h0046};
#218972 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#219372 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0bb, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h1bb, 10'h044, 14'h034b};
#219376 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#219776 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c2, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h220, 10'h044, 14'h0140};
#219780 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#220180 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c8, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h285, 10'h044, 14'h0045};
#220184 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#220584 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ce, 6'h01, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2ea, 10'h044, 14'h014a};
#220588 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#220988 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a2, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02f, 10'h045, 14'h005f};
#220992 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#221392 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a9, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h094, 10'h045, 14'h0054};
#221396 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#221796 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0af, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0f9, 10'h045, 14'h0059};
#221800 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#222200 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0b5, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h15e, 10'h045, 14'h005e};
#222204 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#222604 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0bc, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h1c3, 10'h045, 14'h0353};
#222608 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#223008 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c2, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h228, 10'h045, 14'h0158};
#223012 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#223412 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c8, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h28d, 10'h045, 14'h005d};
#223416 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#223816 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0cf, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2f2, 10'h045, 14'h0052};
#223820 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#224220 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a3, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h037, 10'h046, 14'h0067};
#224224 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#224624 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a9, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h09c, 10'h046, 14'h006c};
#224628 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#225028 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0b0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h101, 10'h046, 14'h0061};
#225032 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#225432 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0b6, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h166, 10'h046, 14'h0366};
#225436 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#225836 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0bc, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h1cb, 10'h046, 14'h036b};
#225840 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#226240 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c3, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h230, 10'h046, 14'h0060};
#226244 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#226644 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c9, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h295, 10'h046, 14'h0065};
#226648 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#227048 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0cf, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2fa, 10'h046, 14'h006a};
#227052 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#227452 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a3, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h03f, 10'h047, 14'h007f};
#227456 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#227856 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0aa, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0a4, 10'h047, 14'h0074};
#227860 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#228260 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0b0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h109, 10'h047, 14'h0079};
#228264 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#228664 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0b6, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h16e, 10'h047, 14'h037e};
#228668 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#229068 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0bd, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1d3, 10'h047, 14'h0073};
#229072 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#229472 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c3, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h238, 10'h047, 14'h0078};
#229476 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#229876 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c9, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h29d, 10'h047, 14'h007d};
#229880 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#230280 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d0, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h302, 10'h047, 14'h0072};
#230284 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#230684 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h047, 10'h048, 14'h0087};
#230688 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#231088 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0aa, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ac, 10'h048, 14'h008c};
#231092 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#231492 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0b1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h111, 10'h048, 14'h0081};
#231496 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#231896 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0b7, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h176, 10'h048, 14'h0386};
#231900 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#232300 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0bd, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1db, 10'h048, 14'h008b};
#232304 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#232704 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h240, 10'h048, 14'h0080};
#232708 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#233108 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ca, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2a5, 10'h048, 14'h0085};
#233112 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#233512 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d0, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h30a, 10'h048, 14'h008a};
#233516 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#233916 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h04f, 10'h049, 14'h009f};
#233920 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#234320 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ab, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0b4, 10'h049, 14'h0094};
#234324 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#234724 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0b1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h119, 10'h049, 14'h0099};
#234728 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#235128 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0b7, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h17e, 10'h049, 14'h039e};
#235132 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#235532 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0be, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1e3, 10'h049, 14'h0093};
#235536 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#235936 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h248, 10'h049, 14'h0098};
#235940 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#236340 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ca, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2ad, 10'h049, 14'h009d};
#236344 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#236744 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d1, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h312, 10'h049, 14'h0092};
#236748 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#237148 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a5, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h057, 10'h04a, 14'h00a7};
#237152 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#237552 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ab, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0bc, 10'h04a, 14'h00ac};
#237556 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#237956 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0b2, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h121, 10'h04a, 14'h02a1};
#237960 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#238360 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0b8, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h186, 10'h04a, 14'h00a6};
#238364 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#238764 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0be, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1eb, 10'h04a, 14'h00ab};
#238768 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#239168 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c5, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h250, 10'h04a, 14'h00a0};
#239172 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#239572 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0cb, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2b5, 10'h04a, 14'h00a5};
#239576 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#239976 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d1, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h31a, 10'h04a, 14'h00aa};
#239980 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#240380 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a5, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h05f, 10'h04b, 14'h00bf};
#240384 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#240784 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ac, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c4, 10'h04b, 14'h00b4};
#240788 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#241188 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0b2, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h129, 10'h04b, 14'h02b9};
#241192 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#241592 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0b8, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h18e, 10'h04b, 14'h00be};
#241596 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#241996 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0bf, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h1f3, 10'h04b, 14'h01b3};
#242000 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#242400 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c5, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h258, 10'h04b, 14'h00b8};
#242404 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#242804 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0cb, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2bd, 10'h04b, 14'h00bd};
#242808 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#243208 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h002, 10'h04c, 14'h00c2};
#243212 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#243612 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a6, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h067, 10'h04c, 14'h00c7};
#243616 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#244016 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ac, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0cc, 10'h04c, 14'h00cc};
#244020 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#244420 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0b3, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h131, 10'h04c, 14'h00c1};
#244424 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#244824 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0b9, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h196, 10'h04c, 14'h00c6};
#244828 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#245228 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0bf, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h1fb, 10'h04c, 14'h01cb};
#245232 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#245632 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c6, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h260, 10'h04c, 14'h00c0};
#245636 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#246036 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0cc, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2c5, 10'h04c, 14'h00c5};
#246040 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#246440 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00a, 10'h04d, 14'h00da};
#246444 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#246844 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a6, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h06f, 10'h04d, 14'h00df};
#246848 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#247248 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ad, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d4, 10'h04d, 14'h00d4};
#247252 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#247652 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0b3, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h139, 10'h04d, 14'h00d9};
#247656 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#248056 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0b9, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h19e, 10'h04d, 14'h00de};
#248060 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#248460 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h203, 10'h04d, 14'h00d3};
#248464 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#248864 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c6, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h268, 10'h04d, 14'h00d8};
#248868 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#249268 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0cc, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2cd, 10'h04d, 14'h00dd};
#249272 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#249672 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h012, 10'h04e, 14'h00e2};
#249676 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#250076 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a7, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h077, 10'h04e, 14'h01e7};
#250080 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#250480 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ad, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0dc, 10'h04e, 14'h00ec};
#250484 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#250884 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0b4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h141, 10'h04e, 14'h00e1};
#250888 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#251288 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ba, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1a6, 10'h04e, 14'h00e6};
#251292 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#251692 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h20b, 10'h04e, 14'h00eb};
#251696 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#252096 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c7, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h270, 10'h04e, 14'h00e0};
#252100 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#252500 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0cd, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2d5, 10'h04e, 14'h00e5};
#252504 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#252904 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h01a, 10'h04f, 14'h00fa};
#252908 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#253308 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0a7, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h07f, 10'h04f, 14'h01ff};
#253312 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#253712 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ae, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h0e4, 10'h04f, 14'h02f4};
#253716 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#254116 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0b4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h149, 10'h04f, 14'h00f9};
#254120 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#254520 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ba, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1ae, 10'h04f, 14'h00fe};
#254524 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#254924 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h213, 10'h04f, 14'h00f3};
#254928 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#255328 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c7, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h278, 10'h04f, 14'h00f8};
#255332 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#255732 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0cd, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2dd, 10'h04f, 14'h00fd};
#255736 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#256136 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ca, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h022, 10'h050, 14'h0002};
#256140 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#256540 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h087, 10'h050, 14'h0007};
#256544 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#256944 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d6, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ec, 10'h050, 14'h000c};
#256948 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#257348 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0dd, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h151, 10'h050, 14'h0001};
#257352 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#257752 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0e3, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1b6, 10'h050, 14'h0006};
#257756 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#258156 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0e9, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h21b, 10'h050, 14'h000b};
#258160 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#258560 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f0, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h280, 10'h050, 14'h0000};
#258564 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#258964 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f6, 6'h01, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2e5, 10'h050, 14'h0105};
#258968 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#259368 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ca, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02a, 10'h051, 14'h001a};
#259372 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#259772 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h08f, 10'h051, 14'h001f};
#259776 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#260176 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d7, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0f4, 10'h051, 14'h0014};
#260180 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#260580 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0dd, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h159, 10'h051, 14'h0019};
#260584 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#260984 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0e3, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1be, 10'h051, 14'h001e};
#260988 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#261388 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ea, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h223, 10'h051, 14'h0113};
#261392 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#261792 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f0, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h288, 10'h051, 14'h0018};
#261796 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#262196 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f6, 6'h01, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2ed, 10'h051, 14'h011d};
#262200 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#262600 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0cb, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h032, 10'h052, 14'h0022};
#262604 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#263004 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h097, 10'h052, 14'h0027};
#263008 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#263408 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d7, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0fc, 10'h052, 14'h002c};
#263412 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#263812 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0de, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h161, 10'h052, 14'h0321};
#263816 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#264216 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0e4, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h1c6, 10'h052, 14'h0326};
#264220 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#264620 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ea, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h22b, 10'h052, 14'h012b};
#264624 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#265024 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f1, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h290, 10'h052, 14'h0020};
#265028 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#265428 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f7, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2f5, 10'h052, 14'h0025};
#265432 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#265832 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0cb, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h03a, 10'h053, 14'h003a};
#265836 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#266236 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h09f, 10'h053, 14'h003f};
#266240 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#266640 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d8, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h104, 10'h053, 14'h0034};
#266644 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#267044 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0de, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h169, 10'h053, 14'h0339};
#267048 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#267448 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0e4, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h1ce, 10'h053, 14'h033e};
#267452 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#267852 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0eb, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h233, 10'h053, 14'h0033};
#267856 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#268256 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f1, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h298, 10'h053, 14'h0038};
#268260 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#268660 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f7, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2fd, 10'h053, 14'h003d};
#268664 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#269064 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0cc, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h042, 10'h054, 14'h0042};
#269068 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#269468 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d2, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0a7, 10'h054, 14'h0047};
#269472 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#269872 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d8, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h10c, 10'h054, 14'h004c};
#269876 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#270276 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0df, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h171, 10'h054, 14'h0041};
#270280 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#270680 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0e5, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1d6, 10'h054, 14'h0046};
#270684 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#271084 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0eb, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h23b, 10'h054, 14'h004b};
#271088 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#271488 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f2, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2a0, 10'h054, 14'h0040};
#271492 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#271892 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f8, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h305, 10'h054, 14'h0045};
#271896 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#272296 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0cc, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h04a, 10'h055, 14'h005a};
#272300 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#272700 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d2, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0af, 10'h055, 14'h005f};
#272704 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#273104 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d9, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h114, 10'h055, 14'h0054};
#273108 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#273508 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0df, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h179, 10'h055, 14'h0059};
#273512 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#273912 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0e5, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1de, 10'h055, 14'h005e};
#273916 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#274316 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ec, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h243, 10'h055, 14'h0053};
#274320 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#274720 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f2, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2a8, 10'h055, 14'h0058};
#274724 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#275124 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f8, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h30d, 10'h055, 14'h005d};
#275128 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#275528 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0cd, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h052, 10'h056, 14'h0062};
#275532 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#275932 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d3, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0b7, 10'h056, 14'h0067};
#275936 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#276336 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d9, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h11c, 10'h056, 14'h006c};
#276340 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#276740 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0e0, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h181, 10'h056, 14'h0361};
#276744 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#277144 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0e6, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1e6, 10'h056, 14'h0066};
#277148 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#277548 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ec, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h24b, 10'h056, 14'h006b};
#277552 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#277952 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f3, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2b0, 10'h056, 14'h0060};
#277956 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#278356 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f9, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h315, 10'h056, 14'h0065};
#278360 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#278760 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0cd, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h05a, 10'h057, 14'h007a};
#278764 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#279164 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d3, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0bf, 10'h057, 14'h007f};
#279168 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#279568 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0da, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h124, 10'h057, 14'h0074};
#279572 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#279972 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0e0, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h189, 10'h057, 14'h0379};
#279976 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#280376 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0e6, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1ee, 10'h057, 14'h007e};
#280380 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#280780 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ed, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h253, 10'h057, 14'h0073};
#280784 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#281184 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f3, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2b8, 10'h057, 14'h0078};
#281188 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#281588 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f9, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h31d, 10'h057, 14'h007d};
#281592 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#281992 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ce, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h062, 10'h058, 14'h0182};
#281996 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#282396 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c7, 10'h058, 14'h0087};
#282400 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#282800 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0da, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h12c, 10'h058, 14'h008c};
#282804 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#283204 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0e1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h191, 10'h058, 14'h0081};
#283208 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#283608 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0e7, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h1f6, 10'h058, 14'h0186};
#283612 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#284012 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ed, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h25b, 10'h058, 14'h008b};
#284016 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#284416 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f4, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2c0, 10'h058, 14'h0080};
#284420 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#284820 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c8, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h005, 10'h059, 14'h0095};
#284824 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#285224 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ce, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h06a, 10'h059, 14'h019a};
#285228 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#285628 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0cf, 10'h059, 14'h009f};
#285632 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#286032 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0db, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h134, 10'h059, 14'h0294};
#286036 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#286436 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0e1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h199, 10'h059, 14'h0099};
#286440 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#286840 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0e7, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h1fe, 10'h059, 14'h019e};
#286844 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#287244 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ee, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h263, 10'h059, 14'h0093};
#287248 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#287648 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f4, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2c8, 10'h059, 14'h0098};
#287652 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#288052 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c8, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00d, 10'h05a, 14'h00ad};
#288056 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#288456 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0cf, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h072, 10'h05a, 14'h00a2};
#288460 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#288860 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d5, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h0d7, 10'h05a, 14'h02a7};
#288864 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#289264 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0db, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h13c, 10'h05a, 14'h02ac};
#289268 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#289668 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0e2, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h1a1, 10'h05a, 14'h03a1};
#289672 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#290072 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0e8, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h206, 10'h05a, 14'h00a6};
#290076 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#290476 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ee, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h26b, 10'h05a, 14'h00ab};
#290480 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#290880 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f5, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2d0, 10'h05a, 14'h00a0};
#290884 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#291284 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c9, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h015, 10'h05b, 14'h00b5};
#291288 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#291688 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0cf, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h07a, 10'h05b, 14'h00ba};
#291692 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#292092 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d5, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h0df, 10'h05b, 14'h02bf};
#292096 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#292496 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0dc, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h144, 10'h05b, 14'h00b4};
#292500 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#292900 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0e2, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h1a9, 10'h05b, 14'h03b9};
#292904 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#293304 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0e8, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h20e, 10'h05b, 14'h00be};
#293308 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#293708 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ef, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h273, 10'h05b, 14'h00b3};
#293712 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#294112 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f5, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2d8, 10'h05b, 14'h00b8};
#294116 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#294516 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0c9, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h01d, 10'h05c, 14'h00cd};
#294520 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#294920 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h082, 10'h05c, 14'h00c2};
#294924 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#295324 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d6, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e7, 10'h05c, 14'h00c7};
#295328 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#295728 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0dc, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h14c, 10'h05c, 14'h00cc};
#295732 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#296132 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0e3, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1b1, 10'h05c, 14'h00c1};
#296136 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#296536 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0e9, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h216, 10'h05c, 14'h00c6};
#296540 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#296940 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ef, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h27b, 10'h05c, 14'h00cb};
#296944 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#297344 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f6, 6'h01, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2e0, 10'h05c, 14'h01c0};
#297348 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#297748 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ca, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h025, 10'h05d, 14'h00d5};
#297752 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#298152 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h08a, 10'h05d, 14'h00da};
#298156 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#298556 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d6, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ef, 10'h05d, 14'h00df};
#298560 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#298960 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0dd, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h154, 10'h05d, 14'h00d4};
#298964 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#299364 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0e3, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1b9, 10'h05d, 14'h00d9};
#299368 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#299768 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0e9, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h21e, 10'h05d, 14'h00de};
#299772 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#300172 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f0, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h283, 10'h05d, 14'h00d3};
#300176 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#300576 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f6, 6'h01, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2e8, 10'h05d, 14'h01d8};
#300580 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#300980 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ca, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02d, 10'h05e, 14'h00ed};
#300984 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#301384 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h092, 10'h05e, 14'h00e2};
#301388 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#301788 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d7, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0f7, 10'h05e, 14'h00e7};
#301792 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#302192 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0dd, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h15c, 10'h05e, 14'h00ec};
#302196 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#302596 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0e4, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h1c1, 10'h05e, 14'h03e1};
#302600 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#303000 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ea, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h226, 10'h05e, 14'h01e6};
#303004 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#303404 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f0, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h28b, 10'h05e, 14'h00eb};
#303408 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#303808 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f7, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2f0, 10'h05e, 14'h00e0};
#303812 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#304212 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0cb, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h035, 10'h05f, 14'h00f5};
#304216 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#304616 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h09a, 10'h05f, 14'h00fa};
#304620 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#305020 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0d7, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ff, 10'h05f, 14'h00ff};
#305024 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#305424 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0de, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h164, 10'h05f, 14'h03f4};
#305428 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#305828 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0e4, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h1c9, 10'h05f, 14'h03f9};
#305832 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#306232 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ea, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h22e, 10'h05f, 14'h01fe};
#306236 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#306636 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f1, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h293, 10'h05f, 14'h00f3};
#306640 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#307040 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f7, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2f8, 10'h05f, 14'h00f8};
#307044 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#307444 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f3, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h03d, 10'h060, 14'h000d};
#307448 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#307848 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0fa, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0a2, 10'h060, 14'h0002};
#307852 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#308252 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h100, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h107, 10'h060, 14'h0007};
#308256 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#308656 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h106, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h16c, 10'h060, 14'h030c};
#308660 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#309060 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h10d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1d1, 10'h060, 14'h0001};
#309064 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#309464 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h113, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h236, 10'h060, 14'h0006};
#309468 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#309868 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h119, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h29b, 10'h060, 14'h000b};
#309872 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#310272 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h120, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h300, 10'h060, 14'h0000};
#310276 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#310676 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h045, 10'h061, 14'h0015};
#310680 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#311080 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0fa, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0aa, 10'h061, 14'h001a};
#311084 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#311484 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h100, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h10f, 10'h061, 14'h001f};
#311488 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#311888 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h107, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h174, 10'h061, 14'h0014};
#311892 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#312292 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h10d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1d9, 10'h061, 14'h0019};
#312296 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#312696 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h113, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h23e, 10'h061, 14'h001e};
#312700 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#313100 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h11a, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2a3, 10'h061, 14'h0013};
#313104 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#313504 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h120, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h308, 10'h061, 14'h0018};
#313508 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#313908 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h04d, 10'h062, 14'h002d};
#313912 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#314312 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0fb, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0b2, 10'h062, 14'h0022};
#314316 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#314716 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h101, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h117, 10'h062, 14'h0027};
#314720 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#315120 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h107, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h17c, 10'h062, 14'h002c};
#315124 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#315524 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h10e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1e1, 10'h062, 14'h0021};
#315528 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#315928 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h114, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h246, 10'h062, 14'h0026};
#315932 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#316332 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h11a, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2ab, 10'h062, 14'h002b};
#316336 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#316736 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h121, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h310, 10'h062, 14'h0020};
#316740 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#317140 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f5, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h055, 10'h063, 14'h0035};
#317144 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#317544 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0fb, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ba, 10'h063, 14'h003a};
#317548 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#317948 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h101, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h11f, 10'h063, 14'h003f};
#317952 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#318352 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h108, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h184, 10'h063, 14'h0034};
#318356 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#318756 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h10e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1e9, 10'h063, 14'h0039};
#318760 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#319160 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h114, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h24e, 10'h063, 14'h003e};
#319164 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#319564 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h11b, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2b3, 10'h063, 14'h0033};
#319568 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#319968 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h121, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h318, 10'h063, 14'h0038};
#319972 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#320372 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f5, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h05d, 10'h064, 14'h004d};
#320376 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#320776 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0fc, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c2, 10'h064, 14'h0042};
#320780 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#321180 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h102, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h127, 10'h064, 14'h0047};
#321184 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#321584 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h108, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h18c, 10'h064, 14'h004c};
#321588 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#321988 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h10f, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h1f1, 10'h064, 14'h0141};
#321992 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#322392 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h115, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h256, 10'h064, 14'h0046};
#322396 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#322796 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h11b, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2bb, 10'h064, 14'h004b};
#322800 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#323200 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h000, 10'h065, 14'h0050};
#323204 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#323604 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f6, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h065, 10'h065, 14'h0155};
#323608 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#324008 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0fc, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ca, 10'h065, 14'h005a};
#324012 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#324412 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h102, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h12f, 10'h065, 14'h005f};
#324416 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#324816 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h109, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h194, 10'h065, 14'h0354};
#324820 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#325220 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h10f, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h1f9, 10'h065, 14'h0159};
#325224 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#325624 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h115, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h25e, 10'h065, 14'h005e};
#325628 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#326028 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h11c, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2c3, 10'h065, 14'h0053};
#326032 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#326432 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h008, 10'h066, 14'h0068};
#326436 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#326836 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f6, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h06d, 10'h066, 14'h016d};
#326840 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#327240 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0fd, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h0d2, 10'h066, 14'h0262};
#327244 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#327644 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h103, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h137, 10'h066, 14'h0267};
#327648 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#328048 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h109, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h19c, 10'h066, 14'h036c};
#328052 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#328452 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h110, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h201, 10'h066, 14'h0161};
#328456 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#328856 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h116, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h266, 10'h066, 14'h0066};
#328860 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#329260 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h11c, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2cb, 10'h066, 14'h006b};
#329264 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#329664 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h010, 10'h067, 14'h0070};
#329668 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#330068 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f7, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h075, 10'h067, 14'h0075};
#330072 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#330472 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0fd, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h0da, 10'h067, 14'h027a};
#330476 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#330876 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h103, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h13f, 10'h067, 14'h027f};
#330880 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#331280 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h10a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1a4, 10'h067, 14'h0074};
#331284 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#331684 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h110, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h209, 10'h067, 14'h0179};
#331688 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#332088 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h116, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h26e, 10'h067, 14'h007e};
#332092 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#332492 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h11d, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2d3, 10'h067, 14'h0073};
#332496 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#332896 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h018, 10'h068, 14'h0088};
#332900 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#333300 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f7, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h07d, 10'h068, 14'h008d};
#333304 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#333704 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0fe, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e2, 10'h068, 14'h0082};
#333708 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#334108 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h104, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h147, 10'h068, 14'h0087};
#334112 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#334512 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h10a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1ac, 10'h068, 14'h008c};
#334516 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#334916 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h111, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h211, 10'h068, 14'h0181};
#334920 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#335320 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h117, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h276, 10'h068, 14'h0086};
#335324 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#335724 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h11d, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2db, 10'h068, 14'h008b};
#335728 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#336128 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f2, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h020, 10'h069, 14'h0090};
#336132 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#336532 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f8, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h085, 10'h069, 14'h0095};
#336536 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#336936 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0fe, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ea, 10'h069, 14'h009a};
#336940 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#337340 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h104, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h14f, 10'h069, 14'h009f};
#337344 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#337744 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h10b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1b4, 10'h069, 14'h0094};
#337748 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#338148 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h111, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h219, 10'h069, 14'h0199};
#338152 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#338552 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h117, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h27e, 10'h069, 14'h009e};
#338556 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#338956 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h11e, 6'h01, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2e3, 10'h069, 14'h0193};
#338960 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#339360 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f2, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h028, 10'h06a, 14'h00a8};
#339364 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#339764 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f8, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h08d, 10'h06a, 14'h00ad};
#339768 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#340168 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ff, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0f2, 10'h06a, 14'h00a2};
#340172 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#340572 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h105, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h157, 10'h06a, 14'h00a7};
#340576 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#340976 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h10b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1bc, 10'h06a, 14'h00ac};
#340980 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#341380 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h112, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h221, 10'h06a, 14'h00a1};
#341384 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#341784 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h118, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h286, 10'h06a, 14'h00a6};
#341788 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#342188 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h11e, 6'h01, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2eb, 10'h06a, 14'h01ab};
#342192 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#342592 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f3, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h030, 10'h06b, 14'h00b0};
#342596 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#342996 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f9, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h095, 10'h06b, 14'h00b5};
#343000 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#343400 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0ff, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0fa, 10'h06b, 14'h00ba};
#343404 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#343804 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h105, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h15f, 10'h06b, 14'h00bf};
#343808 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#344208 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h10c, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h1c4, 10'h06b, 14'h03b4};
#344212 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#344612 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h112, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h229, 10'h06b, 14'h00b9};
#344616 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#345016 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h118, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h28e, 10'h06b, 14'h00be};
#345020 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#345420 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h11f, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2f3, 10'h06b, 14'h00b3};
#345424 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#345824 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f3, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h038, 10'h06c, 14'h00c8};
#345828 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#346228 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f9, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h09d, 10'h06c, 14'h00cd};
#346232 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#346632 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h100, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h102, 10'h06c, 14'h00c2};
#346636 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#347036 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h106, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h167, 10'h06c, 14'h03c7};
#347040 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#347440 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h10c, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h1cc, 10'h06c, 14'h03cc};
#347444 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#347844 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h113, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h231, 10'h06c, 14'h00c1};
#347848 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#348248 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h119, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h296, 10'h06c, 14'h00c6};
#348252 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#348652 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h11f, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2fb, 10'h06c, 14'h00cb};
#348656 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#349056 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h040, 10'h06d, 14'h00d0};
#349060 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#349460 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0fa, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0a5, 10'h06d, 14'h00d5};
#349464 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#349864 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h100, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h10a, 10'h06d, 14'h00da};
#349868 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#350268 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h106, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h16f, 10'h06d, 14'h03df};
#350272 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#350672 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h10d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1d4, 10'h06d, 14'h00d4};
#350676 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#351076 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h113, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h239, 10'h06d, 14'h00d9};
#351080 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#351480 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h119, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h29e, 10'h06d, 14'h00de};
#351484 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#351884 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h120, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h303, 10'h06d, 14'h00d3};
#351888 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#352288 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h048, 10'h06e, 14'h00e8};
#352292 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#352692 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0fa, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ad, 10'h06e, 14'h00ed};
#352696 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#353096 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h101, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h112, 10'h06e, 14'h00e2};
#353100 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#353500 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h107, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h177, 10'h06e, 14'h00e7};
#353504 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#353904 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h10d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1dc, 10'h06e, 14'h00ec};
#353908 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#354308 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h114, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h241, 10'h06e, 14'h00e1};
#354312 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#354712 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h11a, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2a6, 10'h06e, 14'h00e6};
#354716 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#355116 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h120, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h30b, 10'h06e, 14'h00eb};
#355120 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#355520 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0f5, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h050, 10'h06f, 14'h00f0};
#355524 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#355924 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h0fb, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0b5, 10'h06f, 14'h00f5};
#355928 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#356328 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h101, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h11a, 10'h06f, 14'h00fa};
#356332 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#356732 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h107, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h17f, 10'h06f, 14'h00ff};
#356736 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#357136 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h10e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1e4, 10'h06f, 14'h00f4};
#357140 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#357540 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h114, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h249, 10'h06f, 14'h00f9};
#357544 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#357944 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h11a, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2ae, 10'h06f, 14'h00fe};
#357948 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#358348 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h121, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h313, 10'h06f, 14'h00f3};
#358352 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#358752 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h11d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h058, 10'h070, 14'h0008};
#358756 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#359156 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h123, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0bd, 10'h070, 14'h000d};
#359160 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#359560 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h12a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h122, 10'h070, 14'h0002};
#359564 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#359964 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h130, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h187, 10'h070, 14'h0007};
#359968 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#360368 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h136, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1ec, 10'h070, 14'h000c};
#360372 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#360772 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h13d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h251, 10'h070, 14'h0001};
#360776 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#361176 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h143, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2b6, 10'h070, 14'h0006};
#361180 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#361580 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h149, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h31b, 10'h070, 14'h000b};
#361584 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#361984 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h11e, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h060, 10'h071, 14'h0110};
#361988 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#362388 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h124, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c5, 10'h071, 14'h0015};
#362392 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#362792 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h12a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h12a, 10'h071, 14'h001a};
#362796 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#363196 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h130, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h18f, 10'h071, 14'h001f};
#363200 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#363600 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h137, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h1f4, 10'h071, 14'h0114};
#363604 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#364004 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h13d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h259, 10'h071, 14'h0019};
#364008 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#364408 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h143, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2be, 10'h071, 14'h001e};
#364412 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#364812 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h118, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h003, 10'h072, 14'h0023};
#364816 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#365216 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h11e, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h068, 10'h072, 14'h0128};
#365220 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#365620 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h124, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0cd, 10'h072, 14'h002d};
#365624 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#366024 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h12b, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h132, 10'h072, 14'h0222};
#366028 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#366428 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h131, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h197, 10'h072, 14'h0027};
#366432 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#366832 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h137, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h1fc, 10'h072, 14'h012c};
#366836 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#367236 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h13e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h261, 10'h072, 14'h0021};
#367240 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#367640 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h144, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2c6, 10'h072, 14'h0026};
#367644 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#448844 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h14d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d3, 10'h08c, 14'h00c3};
#448848 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#449248 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h153, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h138, 10'h08c, 14'h00c8};
#449252 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#449652 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h159, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h19d, 10'h08c, 14'h00cd};
#449656 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#450056 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h160, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h202, 10'h08c, 14'h00c2};
#450060 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#450460 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h166, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h267, 10'h08c, 14'h00c7};
#450464 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#450864 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h16c, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2cc, 10'h08c, 14'h00cc};
#450868 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#451268 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h141, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h011, 10'h08d, 14'h00d1};
#451272 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#451672 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h147, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h076, 10'h08d, 14'h01d6};
#451676 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#452076 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h14d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0db, 10'h08d, 14'h00db};
#452080 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#452480 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h154, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h140, 10'h08d, 14'h00d0};
#452484 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#452884 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h15a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1a5, 10'h08d, 14'h00d5};
#452888 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#453288 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h160, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h20a, 10'h08d, 14'h00da};
#453292 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#453692 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h166, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h26f, 10'h08d, 14'h00df};
#453696 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#454096 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h16d, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2d4, 10'h08d, 14'h00d4};
#454100 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#454500 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h141, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h019, 10'h08e, 14'h00e9};
#454504 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#454904 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h147, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h07e, 10'h08e, 14'h01ee};
#454908 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#455308 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h14e, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h0e3, 10'h08e, 14'h02e3};
#455312 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#455712 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h154, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h148, 10'h08e, 14'h00e8};
#455716 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#456116 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h15a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1ad, 10'h08e, 14'h00ed};
#456120 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#456520 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h161, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h212, 10'h08e, 14'h00e2};
#456524 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#456924 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h167, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h277, 10'h08e, 14'h00e7};
#456928 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#457328 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h16d, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2dc, 10'h08e, 14'h00ec};
#457332 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#457732 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h142, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h021, 10'h08f, 14'h00f1};
#457736 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#458136 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h148, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h086, 10'h08f, 14'h00f6};
#458140 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#458540 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h14e, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h0eb, 10'h08f, 14'h02fb};
#458544 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#458944 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h155, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h150, 10'h08f, 14'h00f0};
#458948 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#459348 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h15b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1b5, 10'h08f, 14'h00f5};
#459352 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#459752 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h161, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h21a, 10'h08f, 14'h00fa};
#459756 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#460156 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h167, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h27f, 10'h08f, 14'h00ff};
#460160 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#460560 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h16e, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2e4, 10'h08f, 14'h00f4};
#460564 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#460964 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h16a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h029, 10'h090, 14'h0009};
#460968 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#461368 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h170, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h08e, 10'h090, 14'h010e};
#461372 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#461772 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h177, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h0f3, 10'h090, 14'h0203};
#461776 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#462176 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h17d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h158, 10'h090, 14'h0008};
#462180 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#462580 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h183, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1bd, 10'h090, 14'h000d};
#462584 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#462984 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h18a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h222, 10'h090, 14'h0002};
#462988 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#463388 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h190, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h287, 10'h090, 14'h0007};
#463392 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#463792 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h196, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2ec, 10'h090, 14'h000c};
#463796 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#464196 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h16b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h031, 10'h091, 14'h0011};
#464200 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#464600 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h171, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h096, 10'h091, 14'h0116};
#464604 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#465004 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h177, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h0fb, 10'h091, 14'h021b};
#465008 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#465408 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h17e, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h160, 10'h091, 14'h0310};
#465412 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#465812 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h184, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h1c5, 10'h091, 14'h0315};
#465816 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#466216 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h18a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h22a, 10'h091, 14'h001a};
#466220 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#466620 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h190, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h28f, 10'h091, 14'h001f};
#466624 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#467024 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h197, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2f4, 10'h091, 14'h0014};
#467028 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#467428 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h16b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h039, 10'h092, 14'h0029};
#467432 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#467832 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h171, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h09e, 10'h092, 14'h012e};
#467836 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#468236 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h178, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h103, 10'h092, 14'h0223};
#468240 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#468640 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h17e, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h168, 10'h092, 14'h0328};
#468644 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#549844 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1b9, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h295, 10'h0ab, 14'h00b5};
#549848 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#550248 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1bf, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2fa, 10'h0ab, 14'h00ba};
#550252 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#550652 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h193, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h03f, 10'h0ac, 14'h00cf};
#550656 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#551056 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h19a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0a4, 10'h0ac, 14'h00c4};
#551060 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#551460 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1a0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h109, 10'h0ac, 14'h00c9};
#551464 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#551864 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1a6, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h16e, 10'h0ac, 14'h00ce};
#551868 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#552268 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1ad, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1d3, 10'h0ac, 14'h00c3};
#552272 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#552672 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1b3, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h238, 10'h0ac, 14'h00c8};
#552676 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#553076 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1b9, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h29d, 10'h0ac, 14'h00cd};
#553080 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#553480 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1c0, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h302, 10'h0ac, 14'h00c2};
#553484 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#553884 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h194, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h047, 10'h0ad, 14'h00d7};
#553888 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#554288 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h19a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ac, 10'h0ad, 14'h00dc};
#554292 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#554692 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1a1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h111, 10'h0ad, 14'h00d1};
#554696 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#555096 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1a7, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h176, 10'h0ad, 14'h00d6};
#555100 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#555500 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1ad, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1db, 10'h0ad, 14'h00db};
#555504 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#555904 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1b4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h240, 10'h0ad, 14'h00d0};
#555908 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#556308 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1ba, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2a5, 10'h0ad, 14'h00d5};
#556312 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#556712 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1c0, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h30a, 10'h0ad, 14'h00da};
#556716 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#557116 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h194, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h04f, 10'h0ae, 14'h00ef};
#557120 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#557520 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h19b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0b4, 10'h0ae, 14'h00e4};
#557524 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#557924 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1a1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h119, 10'h0ae, 14'h00e9};
#557928 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#558328 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1a7, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h17e, 10'h0ae, 14'h00ee};
#558332 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#558732 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1ae, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1e3, 10'h0ae, 14'h00e3};
#558736 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#559136 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1b4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h248, 10'h0ae, 14'h00e8};
#559140 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#559540 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1ba, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2ad, 10'h0ae, 14'h00ed};
#559544 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#559944 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1c1, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h312, 10'h0ae, 14'h00e2};
#559948 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#560348 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h195, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h057, 10'h0af, 14'h00f7};
#560352 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#560752 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h19b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0bc, 10'h0af, 14'h00fc};
#560756 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#561156 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1a2, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h121, 10'h0af, 14'h00f1};
#561160 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#561560 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1a8, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h186, 10'h0af, 14'h00f6};
#561564 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#561964 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1ae, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1eb, 10'h0af, 14'h00fb};
#561968 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#562368 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1b5, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h250, 10'h0af, 14'h00f0};
#562372 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#562772 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1bb, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2b5, 10'h0af, 14'h00f5};
#562776 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#563176 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1c1, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h31a, 10'h0af, 14'h00fa};
#563180 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#563580 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1bd, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h05f, 10'h0b0, 14'h000f};
#563584 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#563984 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1c4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c4, 10'h0b0, 14'h0004};
#563988 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#564388 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1ca, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h129, 10'h0b0, 14'h0009};
#564392 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#564792 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1d0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h18e, 10'h0b0, 14'h000e};
#564796 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#565196 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1d7, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1f3, 10'h0b0, 14'h0003};
#565200 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#565600 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1dd, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h258, 10'h0b0, 14'h0008};
#565604 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#566004 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1e3, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2bd, 10'h0b0, 14'h000d};
#566008 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#566408 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1b8, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h002, 10'h0b1, 14'h0012};
#566412 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#566812 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1be, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h067, 10'h0b1, 14'h0017};
#566816 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#567216 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1c4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0cc, 10'h0b1, 14'h001c};
#567220 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#567620 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1cb, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h131, 10'h0b1, 14'h0011};
#567624 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#568024 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1d1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h196, 10'h0b1, 14'h0016};
#568028 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#568428 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1d7, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1fb, 10'h0b1, 14'h001b};
#568432 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#568832 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1de, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h260, 10'h0b1, 14'h0010};
#568836 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#569236 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1e4, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2c5, 10'h0b1, 14'h0015};
#569240 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#569640 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1b8, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00a, 10'h0b2, 14'h002a};
#569644 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#650844 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1f3, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h137, 10'h0cb, 14'h00b7};
#650848 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#651248 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1f9, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h19c, 10'h0cb, 14'h00bc};
#651252 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#651652 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h200, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h201, 10'h0cb, 14'h00b1};
#651656 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#652056 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h206, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h266, 10'h0cb, 14'h00b6};
#652060 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#652460 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h20c, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2cb, 10'h0cb, 14'h00bb};
#652464 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#652864 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1e1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h010, 10'h0cc, 14'h00c0};
#652868 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#653268 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1e7, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h075, 10'h0cc, 14'h00c5};
#653272 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#653672 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1ed, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0da, 10'h0cc, 14'h00ca};
#653676 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#654076 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1f3, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h13f, 10'h0cc, 14'h00cf};
#654080 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#654480 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1fa, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1a4, 10'h0cc, 14'h00c4};
#654484 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#654884 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h200, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h209, 10'h0cc, 14'h00c9};
#654888 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#655288 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h206, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h26e, 10'h0cc, 14'h00ce};
#655292 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#655692 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h20d, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2d3, 10'h0cc, 14'h00c3};
#655696 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#656096 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1e1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h018, 10'h0cd, 14'h00d8};
#656100 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#656500 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1e7, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h07d, 10'h0cd, 14'h00dd};
#656504 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#656904 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1ee, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e2, 10'h0cd, 14'h00d2};
#656908 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#657308 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1f4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h147, 10'h0cd, 14'h00d7};
#657312 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#657712 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1fa, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1ac, 10'h0cd, 14'h00dc};
#657716 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#658116 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h201, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h211, 10'h0cd, 14'h00d1};
#658120 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#658520 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h207, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h276, 10'h0cd, 14'h00d6};
#658524 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#658924 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h20d, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2db, 10'h0cd, 14'h00db};
#658928 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#659328 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1e2, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h020, 10'h0ce, 14'h00e0};
#659332 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#659732 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1e8, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h085, 10'h0ce, 14'h00e5};
#659736 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#660136 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1ee, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ea, 10'h0ce, 14'h00ea};
#660140 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#660540 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1f4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h14f, 10'h0ce, 14'h00ef};
#660544 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#660944 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1fb, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1b4, 10'h0ce, 14'h00e4};
#660948 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#661348 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h201, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h219, 10'h0ce, 14'h00e9};
#661352 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#661752 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h207, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h27e, 10'h0ce, 14'h00ee};
#661756 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#662156 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h20e, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2e3, 10'h0ce, 14'h00e3};
#662160 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#662560 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1e2, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h028, 10'h0cf, 14'h00f8};
#662564 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#662964 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1e8, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h08d, 10'h0cf, 14'h00fd};
#662968 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#663368 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1ef, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0f2, 10'h0cf, 14'h00f2};
#663372 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#663772 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1f5, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h157, 10'h0cf, 14'h00f7};
#663776 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#664176 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h1fb, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1bc, 10'h0cf, 14'h00fc};
#664180 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#664580 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h202, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h221, 10'h0cf, 14'h00f1};
#664584 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#664984 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h208, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h286, 10'h0cf, 14'h00f6};
#664988 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#665388 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h20e, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2eb, 10'h0cf, 14'h00fb};
#665392 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#665792 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h20b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h030, 10'h0d0, 14'h0000};
#665796 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#666196 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h211, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h095, 10'h0d0, 14'h0005};
#666200 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#666600 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h217, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h0fa, 10'h0d0, 14'h020a};
#666604 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#667004 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h21d, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h15f, 10'h0d0, 14'h030f};
#667008 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#667408 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h224, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1c4, 10'h0d0, 14'h0004};
#667412 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#667812 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h22a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h229, 10'h0d0, 14'h0009};
#667816 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#668216 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h230, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h28e, 10'h0d0, 14'h000e};
#668220 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#668620 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h237, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2f3, 10'h0d0, 14'h0003};
#668624 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#669024 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h20b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h038, 10'h0d1, 14'h0018};
#669028 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#669428 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h211, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h09d, 10'h0d1, 14'h001d};
#669432 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#669832 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h218, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h102, 10'h0d1, 14'h0012};
#669836 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#670236 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h21e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h167, 10'h0d1, 14'h0017};
#670240 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#670640 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h224, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1cc, 10'h0d1, 14'h001c};
#670644 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#751844 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h25f, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2f9, 10'h0ea, 14'h00a9};
#751848 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#752248 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h233, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h03e, 10'h0eb, 14'h00be};
#752252 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#752652 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h23a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0a3, 10'h0eb, 14'h00b3};
#752656 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#753056 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h240, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h108, 10'h0eb, 14'h00b8};
#753060 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#753460 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h246, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h16d, 10'h0eb, 14'h00bd};
#753464 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#753864 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h24d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1d2, 10'h0eb, 14'h00b2};
#753868 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#754268 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h253, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h237, 10'h0eb, 14'h00b7};
#754272 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#754672 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h259, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h29c, 10'h0eb, 14'h00bc};
#754676 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#755076 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h260, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h301, 10'h0eb, 14'h00b1};
#755080 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#755480 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h234, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h046, 10'h0ec, 14'h00c6};
#755484 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#755884 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h23a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ab, 10'h0ec, 14'h00cb};
#755888 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#756288 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h241, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h110, 10'h0ec, 14'h00c0};
#756292 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#756692 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h247, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h175, 10'h0ec, 14'h00c5};
#756696 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#757096 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h24d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1da, 10'h0ec, 14'h00ca};
#757100 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#757500 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h253, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h23f, 10'h0ec, 14'h00cf};
#757504 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#757904 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h25a, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2a4, 10'h0ec, 14'h00c4};
#757908 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#758308 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h260, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h309, 10'h0ec, 14'h00c9};
#758312 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#758712 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h234, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h04e, 10'h0ed, 14'h00de};
#758716 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#759116 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h23b, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h0b3, 10'h0ed, 14'h02d3};
#759120 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#759520 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h241, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h118, 10'h0ed, 14'h00d8};
#759524 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#759924 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h247, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h17d, 10'h0ed, 14'h00dd};
#759928 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#760328 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h24e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1e2, 10'h0ed, 14'h00d2};
#760332 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#760732 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h254, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h247, 10'h0ed, 14'h00d7};
#760736 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#761136 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h25a, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2ac, 10'h0ed, 14'h00dc};
#761140 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#761540 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h261, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h311, 10'h0ed, 14'h00d1};
#761544 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#761944 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h235, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h056, 10'h0ee, 14'h00e6};
#761948 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#762348 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h23b, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h0bb, 10'h0ee, 14'h02eb};
#762352 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#762752 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h242, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h120, 10'h0ee, 14'h00e0};
#762756 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#763156 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h248, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h185, 10'h0ee, 14'h00e5};
#763160 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#763560 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h24e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1ea, 10'h0ee, 14'h00ea};
#763564 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#763964 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h254, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h24f, 10'h0ee, 14'h00ef};
#763968 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#764368 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h25b, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2b4, 10'h0ee, 14'h00e4};
#764372 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#764772 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h261, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h319, 10'h0ee, 14'h00e9};
#764776 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#765176 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h235, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h05e, 10'h0ef, 14'h00fe};
#765180 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#765580 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h23c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c3, 10'h0ef, 14'h00f3};
#765584 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#765984 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h242, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h128, 10'h0ef, 14'h00f8};
#765988 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#766388 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h248, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h18d, 10'h0ef, 14'h00fd};
#766392 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#766792 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h24f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1f2, 10'h0ef, 14'h00f2};
#766796 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#767196 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h255, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h257, 10'h0ef, 14'h00f7};
#767200 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#767600 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h25b, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2bc, 10'h0ef, 14'h00fc};
#767604 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#768004 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h258, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h001, 10'h0f0, 14'h0001};
#768008 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#768408 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h25e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h066, 10'h0f0, 14'h0006};
#768412 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#768812 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h264, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h0cb, 10'h0f0, 14'h020b};
#768816 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#769216 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h26b, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h130, 10'h0f0, 14'h0300};
#769220 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#769620 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h271, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h195, 10'h0f0, 14'h0005};
#769624 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#770024 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h277, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1fa, 10'h0f0, 14'h000a};
#770028 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#770428 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h27d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h25f, 10'h0f0, 14'h000f};
#770432 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#770832 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h284, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2c4, 10'h0f0, 14'h0004};
#770836 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#771236 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h258, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h009, 10'h0f1, 14'h0019};
#771240 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#771640 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h25e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h06e, 10'h0f1, 14'h001e};
#771644 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#852844 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h299, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h19b, 10'h10a, 14'h00ab};
#852848 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#853248 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2a0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h200, 10'h10a, 14'h00a0};
#853252 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#853652 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2a6, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h265, 10'h10a, 14'h00a5};
#853656 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#854056 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2ac, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2ca, 10'h10a, 14'h00aa};
#854060 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#854460 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h280, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00f, 10'h10b, 14'h00bf};
#854464 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#854864 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h287, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h074, 10'h10b, 14'h00b4};
#854868 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#855268 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h28d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d9, 10'h10b, 14'h00b9};
#855272 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#855672 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h293, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h13e, 10'h10b, 14'h00be};
#855676 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#856076 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h29a, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h1a3, 10'h10b, 14'h01b3};
#856080 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#856480 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2a0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h208, 10'h10b, 14'h00b8};
#856484 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#856884 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2a6, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h26d, 10'h10b, 14'h00bd};
#856888 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#857288 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2ad, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2d2, 10'h10b, 14'h00b2};
#857292 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#857692 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h281, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h017, 10'h10c, 14'h00c7};
#857696 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#858096 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h287, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h07c, 10'h10c, 14'h00cc};
#858100 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#858500 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h28e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e1, 10'h10c, 14'h00c1};
#858504 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#858904 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h294, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h146, 10'h10c, 14'h00c6};
#858908 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#859308 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h29a, 6'h01, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h1ab, 10'h10c, 14'h01cb};
#859312 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#859712 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2a1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h210, 10'h10c, 14'h00c0};
#859716 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#860116 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2a7, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h275, 10'h10c, 14'h00c5};
#860120 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#860520 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2ad, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2da, 10'h10c, 14'h00ca};
#860524 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#860924 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h281, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h01f, 10'h10d, 14'h00df};
#860928 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#861328 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h288, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h084, 10'h10d, 14'h00d4};
#861332 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#861732 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h28e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e9, 10'h10d, 14'h00d9};
#861736 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#862136 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h294, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h14e, 10'h10d, 14'h00de};
#862140 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#862540 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h29b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1b3, 10'h10d, 14'h00d3};
#862544 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#862944 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2a1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h218, 10'h10d, 14'h00d8};
#862948 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#863348 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2a7, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h27d, 10'h10d, 14'h00dd};
#863352 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#863752 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2ae, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2e2, 10'h10d, 14'h00d2};
#863756 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#864156 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h282, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h027, 10'h10e, 14'h00e7};
#864160 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#864560 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h288, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h08c, 10'h10e, 14'h00ec};
#864564 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#864964 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h28f, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h0f1, 10'h10e, 14'h02e1};
#864968 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#865368 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h295, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h156, 10'h10e, 14'h03e6};
#865372 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#865772 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h29b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1bb, 10'h10e, 14'h00eb};
#865776 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#866176 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2a2, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h220, 10'h10e, 14'h00e0};
#866180 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#866580 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2a8, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h285, 10'h10e, 14'h00e5};
#866584 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#866984 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2ae, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2ea, 10'h10e, 14'h00ea};
#866988 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#867388 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h282, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02f, 10'h10f, 14'h00ff};
#867392 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#867792 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h289, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h094, 10'h10f, 14'h00f4};
#867796 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#868196 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h28f, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h0f9, 10'h10f, 14'h02f9};
#868200 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#868600 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h295, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h15e, 10'h10f, 14'h03fe};
#868604 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#869004 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h29c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1c3, 10'h10f, 14'h00f3};
#869008 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#869408 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2a2, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h228, 10'h10f, 14'h00f8};
#869412 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#869812 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2a8, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h28d, 10'h10f, 14'h00fd};
#869816 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#870216 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2af, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2f2, 10'h10f, 14'h00f2};
#870220 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#870620 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2ab, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h037, 10'h110, 14'h0007};
#870624 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#871024 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2b1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h09c, 10'h110, 14'h000c};
#871028 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#871428 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2b8, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h101, 10'h110, 14'h0001};
#871432 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#871832 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2be, 6'h03, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h166, 10'h110, 14'h0306};
#871836 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#872236 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2c4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1cb, 10'h110, 14'h000b};
#872240 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#872640 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2cb, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h230, 10'h110, 14'h0000};
#872644 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#953844 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2d3, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h03d, 10'h12a, 14'h00ad};
#953848 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#954248 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2da, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0a2, 10'h12a, 14'h00a2};
#954252 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#954652 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2e0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h107, 10'h12a, 14'h00a7};
#954656 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#955056 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2e6, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h16c, 10'h12a, 14'h00ac};
#955060 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#955460 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2ed, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1d1, 10'h12a, 14'h00a1};
#955464 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#955864 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2f3, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h236, 10'h12a, 14'h00a6};
#955868 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#956268 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2f9, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h29b, 10'h12a, 14'h00ab};
#956272 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#956672 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h300, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h300, 10'h12a, 14'h00a0};
#956676 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#957076 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2d4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h045, 10'h12b, 14'h00b5};
#957080 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#957480 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2da, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0aa, 10'h12b, 14'h00ba};
#957484 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#957884 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2e0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h10f, 10'h12b, 14'h00bf};
#957888 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#958288 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2e7, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h174, 10'h12b, 14'h00b4};
#958292 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#958692 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2ed, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1d9, 10'h12b, 14'h00b9};
#958696 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#959096 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2f3, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h23e, 10'h12b, 14'h00be};
#959100 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#959500 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2fa, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2a3, 10'h12b, 14'h00b3};
#959504 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#959904 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h300, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h308, 10'h12b, 14'h00b8};
#959908 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#960308 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2d4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h04d, 10'h12c, 14'h00cd};
#960312 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#960712 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2db, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h0b2, 10'h12c, 14'h02c2};
#960716 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#961116 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2e1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h117, 10'h12c, 14'h00c7};
#961120 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#961520 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2e7, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h17c, 10'h12c, 14'h00cc};
#961524 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#961924 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2ee, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1e1, 10'h12c, 14'h00c1};
#961928 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#962328 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2f4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h246, 10'h12c, 14'h00c6};
#962332 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#962732 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2fa, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2ab, 10'h12c, 14'h00cb};
#962736 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#963136 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h301, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h310, 10'h12c, 14'h00c0};
#963140 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#963540 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2d5, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h055, 10'h12d, 14'h00d5};
#963544 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#963944 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2db, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h0ba, 10'h12d, 14'h02da};
#963948 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#964348 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2e1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h11f, 10'h12d, 14'h00df};
#964352 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#964752 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2e8, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h184, 10'h12d, 14'h00d4};
#964756 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#965156 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2ee, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1e9, 10'h12d, 14'h00d9};
#965160 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#965560 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2f4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h24e, 10'h12d, 14'h00de};
#965564 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#965964 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2fb, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2b3, 10'h12d, 14'h00d3};
#965968 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#966368 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h301, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h318, 10'h12d, 14'h00d8};
#966372 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#966772 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2d5, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h05d, 10'h12e, 14'h00ed};
#966776 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#967176 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2dc, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c2, 10'h12e, 14'h00e2};
#967180 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#967580 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2e2, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h127, 10'h12e, 14'h00e7};
#967584 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#967984 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2e8, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h18c, 10'h12e, 14'h00ec};
#967988 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#968388 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2ef, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1f1, 10'h12e, 14'h00e1};
#968392 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#968792 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2f5, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h256, 10'h12e, 14'h00e6};
#968796 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#969196 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2fb, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2bb, 10'h12e, 14'h00eb};
#969200 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#969600 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2d0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h000, 10'h12f, 14'h00f0};
#969604 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#970004 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2d6, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h065, 10'h12f, 14'h00f5};
#970008 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#970408 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2dc, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ca, 10'h12f, 14'h00fa};
#970412 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#970812 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2e2, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h12f, 10'h12f, 14'h00ff};
#970816 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#971216 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2e9, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h194, 10'h12f, 14'h00f4};
#971220 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#971620 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2ef, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1f9, 10'h12f, 14'h00f9};
#971624 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#972024 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2f5, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h25e, 10'h12f, 14'h00fe};
#972028 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#972428 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2fc, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2c3, 10'h12f, 14'h00f3};
#972432 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#972832 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2f8, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h008, 10'h130, 14'h0008};
#972836 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#973236 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h2fe, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h06d, 10'h130, 14'h000d};
#973240 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#973640 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h305, 6'h02, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h0d2, 10'h130, 14'h0202};
#973644 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1054844 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h33f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1ff, 10'h149, 14'h009f};
#1054848 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1055248 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h346, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h264, 10'h149, 14'h0094};
#1055252 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1055652 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h34c, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2c9, 10'h149, 14'h0099};
#1055656 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1056056 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h320, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00e, 10'h14a, 14'h00ae};
#1056060 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1056460 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h327, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h073, 10'h14a, 14'h00a3};
#1056464 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1056864 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h32d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d8, 10'h14a, 14'h00a8};
#1056868 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1057268 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h333, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h13d, 10'h14a, 14'h00ad};
#1057272 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1057672 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h33a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1a2, 10'h14a, 14'h00a2};
#1057676 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1058076 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h340, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h207, 10'h14a, 14'h00a7};
#1058080 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1058480 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h346, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h26c, 10'h14a, 14'h00ac};
#1058484 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1058884 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h34d, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2d1, 10'h14a, 14'h00a1};
#1058888 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1059288 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h321, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h016, 10'h14b, 14'h00b6};
#1059292 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1059692 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h327, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h07b, 10'h14b, 14'h00bb};
#1059696 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1060096 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h32e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e0, 10'h14b, 14'h00b0};
#1060100 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1060500 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h334, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h145, 10'h14b, 14'h00b5};
#1060504 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1060904 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h33a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1aa, 10'h14b, 14'h00ba};
#1060908 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1061308 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h340, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h20f, 10'h14b, 14'h00bf};
#1061312 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1061712 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h347, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h274, 10'h14b, 14'h00b4};
#1061716 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1062116 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h34d, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2d9, 10'h14b, 14'h00b9};
#1062120 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1062520 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h321, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h01e, 10'h14c, 14'h00ce};
#1062524 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1062924 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h328, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h083, 10'h14c, 14'h00c3};
#1062928 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1063328 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h32e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e8, 10'h14c, 14'h00c8};
#1063332 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1063732 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h334, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h14d, 10'h14c, 14'h00cd};
#1063736 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1064136 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h33b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1b2, 10'h14c, 14'h00c2};
#1064140 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1064540 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h341, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h217, 10'h14c, 14'h00c7};
#1064544 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1064944 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h347, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h27c, 10'h14c, 14'h00cc};
#1064948 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1065348 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h34e, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2e1, 10'h14c, 14'h00c1};
#1065352 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1065752 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h322, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h026, 10'h14d, 14'h00d6};
#1065756 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1066156 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h328, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h08b, 10'h14d, 14'h00db};
#1066160 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1066560 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h32f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0f0, 10'h14d, 14'h00d0};
#1066564 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1066964 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h335, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h155, 10'h14d, 14'h00d5};
#1066968 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1067368 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h33b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1ba, 10'h14d, 14'h00da};
#1067372 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1067772 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h341, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h21f, 10'h14d, 14'h00df};
#1067776 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1068176 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h348, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h284, 10'h14d, 14'h00d4};
#1068180 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1068580 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h34e, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2e9, 10'h14d, 14'h00d9};
#1068584 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1068984 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h322, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02e, 10'h14e, 14'h00ee};
#1068988 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1069388 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h329, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h093, 10'h14e, 14'h00e3};
#1069392 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1069792 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h32f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0f8, 10'h14e, 14'h00e8};
#1069796 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1070196 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h335, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h15d, 10'h14e, 14'h00ed};
#1070200 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1070600 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h33c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1c2, 10'h14e, 14'h00e2};
#1070604 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1071004 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h342, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h227, 10'h14e, 14'h00e7};
#1071008 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1071408 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h348, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h28c, 10'h14e, 14'h00ec};
#1071412 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1071812 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h34f, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2f1, 10'h14e, 14'h00e1};
#1071816 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1072216 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h323, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h036, 10'h14f, 14'h00f6};
#1072220 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1072620 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h329, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h09b, 10'h14f, 14'h00fb};
#1072624 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1073024 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h330, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h100, 10'h14f, 14'h00f0};
#1073028 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1073428 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h336, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h165, 10'h14f, 14'h00f5};
#1073432 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1073832 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h33c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1ca, 10'h14f, 14'h00fa};
#1073836 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1074236 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h342, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h22f, 10'h14f, 14'h00ff};
#1074240 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1074640 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h349, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h294, 10'h14f, 14'h00f4};
#1074644 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1155844 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h37a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0a1, 10'h169, 14'h0091};
#1155848 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1156248 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h380, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h106, 10'h169, 14'h0096};
#1156252 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1156652 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h386, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h16b, 10'h169, 14'h009b};
#1156656 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1157056 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h38d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1d0, 10'h169, 14'h0090};
#1157060 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1157460 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h393, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h235, 10'h169, 14'h0095};
#1157464 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1157864 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h399, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h29a, 10'h169, 14'h009a};
#1157868 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1158268 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h39f, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2ff, 10'h169, 14'h009f};
#1158272 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1158672 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h374, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h044, 10'h16a, 14'h00a4};
#1158676 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1159076 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h37a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0a9, 10'h16a, 14'h00a9};
#1159080 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1159480 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h380, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h10e, 10'h16a, 14'h00ae};
#1159484 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1159884 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h387, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h173, 10'h16a, 14'h00a3};
#1159888 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1160288 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h38d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1d8, 10'h16a, 14'h00a8};
#1160292 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1160692 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h393, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h23d, 10'h16a, 14'h00ad};
#1160696 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1161096 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h39a, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2a2, 10'h16a, 14'h00a2};
#1161100 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1161500 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3a0, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h307, 10'h16a, 14'h00a7};
#1161504 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1161904 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h374, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h04c, 10'h16b, 14'h00bc};
#1161908 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1162308 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h37b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0b1, 10'h16b, 14'h00b1};
#1162312 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1162712 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h381, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h116, 10'h16b, 14'h00b6};
#1162716 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1163116 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h387, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h17b, 10'h16b, 14'h00bb};
#1163120 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1163520 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h38e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1e0, 10'h16b, 14'h00b0};
#1163524 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1163924 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h394, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h245, 10'h16b, 14'h00b5};
#1163928 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1164328 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h39a, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2aa, 10'h16b, 14'h00ba};
#1164332 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1164732 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3a0, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h30f, 10'h16b, 14'h00bf};
#1164736 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1165136 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h375, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h054, 10'h16c, 14'h00c4};
#1165140 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1165540 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h37b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0b9, 10'h16c, 14'h00c9};
#1165544 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1165944 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h381, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h11e, 10'h16c, 14'h00ce};
#1165948 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1166348 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h388, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h183, 10'h16c, 14'h00c3};
#1166352 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1166752 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h38e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1e8, 10'h16c, 14'h00c8};
#1166756 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1167156 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h394, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h24d, 10'h16c, 14'h00cd};
#1167160 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1167560 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h39b, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2b2, 10'h16c, 14'h00c2};
#1167564 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1167964 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3a1, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h317, 10'h16c, 14'h00c7};
#1167968 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1168368 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h375, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h05c, 10'h16d, 14'h00dc};
#1168372 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1168772 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h37c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c1, 10'h16d, 14'h00d1};
#1168776 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1169176 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h382, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h126, 10'h16d, 14'h00d6};
#1169180 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1169580 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h388, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h18b, 10'h16d, 14'h00db};
#1169584 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1169984 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h38f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1f0, 10'h16d, 14'h00d0};
#1169988 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1170388 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h395, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h255, 10'h16d, 14'h00d5};
#1170392 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1170792 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h39b, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2ba, 10'h16d, 14'h00da};
#1170796 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1171196 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3a1, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h31f, 10'h16d, 14'h00df};
#1171200 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1171600 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h376, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h064, 10'h16e, 14'h00e4};
#1171604 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1172004 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h37c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c9, 10'h16e, 14'h00e9};
#1172008 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1172408 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h382, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h12e, 10'h16e, 14'h00ee};
#1172412 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1172812 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h389, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h193, 10'h16e, 14'h00e3};
#1172816 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1173216 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h38f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1f8, 10'h16e, 14'h00e8};
#1173220 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1173620 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h395, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h25d, 10'h16e, 14'h00ed};
#1173624 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1174024 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h39c, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2c2, 10'h16e, 14'h00e2};
#1174028 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1174428 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h370, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h007, 10'h16f, 14'h00f7};
#1174432 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1174832 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h376, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h06c, 10'h16f, 14'h00fc};
#1174836 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1175236 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h37d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d1, 10'h16f, 14'h00f1};
#1175240 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1175640 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h383, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h136, 10'h16f, 14'h00f6};
#1175644 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1256844 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3e6, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h263, 10'h188, 14'h0083};
#1256848 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1257248 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3ec, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2c8, 10'h188, 14'h0088};
#1257252 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1257652 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3c0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00d, 10'h189, 14'h009d};
#1257656 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1258056 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3c7, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h072, 10'h189, 14'h0092};
#1258060 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1258460 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3cd, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d7, 10'h189, 14'h0097};
#1258464 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1258864 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3d3, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h13c, 10'h189, 14'h009c};
#1258868 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1259268 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3da, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1a1, 10'h189, 14'h0091};
#1259272 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1259672 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3e0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h206, 10'h189, 14'h0096};
#1259676 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1260076 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3e6, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h26b, 10'h189, 14'h009b};
#1260080 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1260480 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3ed, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2d0, 10'h189, 14'h0090};
#1260484 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1260884 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3c1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h015, 10'h18a, 14'h00a5};
#1260888 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1261288 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3c7, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h07a, 10'h18a, 14'h00aa};
#1261292 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1261692 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3cd, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0df, 10'h18a, 14'h00af};
#1261696 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1262096 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3d4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h144, 10'h18a, 14'h00a4};
#1262100 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1262500 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3da, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1a9, 10'h18a, 14'h00a9};
#1262504 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1262904 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3e0, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h20e, 10'h18a, 14'h00ae};
#1262908 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1263308 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3e7, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h273, 10'h18a, 14'h00a3};
#1263312 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1263712 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3ed, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2d8, 10'h18a, 14'h00a8};
#1263716 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1264116 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3c1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h01d, 10'h18b, 14'h00bd};
#1264120 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1264520 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3c8, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h082, 10'h18b, 14'h00b2};
#1264524 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1264924 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3ce, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e7, 10'h18b, 14'h00b7};
#1264928 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1265328 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3d4, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h14c, 10'h18b, 14'h00bc};
#1265332 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1265732 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3db, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1b1, 10'h18b, 14'h00b1};
#1265736 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1266136 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3e1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h216, 10'h18b, 14'h00b6};
#1266140 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1266540 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3e7, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h27b, 10'h18b, 14'h00bb};
#1266544 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1266944 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3ee, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2e0, 10'h18b, 14'h00b0};
#1266948 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1267348 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3c2, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h025, 10'h18c, 14'h00c5};
#1267352 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1267752 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3c8, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h08a, 10'h18c, 14'h00ca};
#1267756 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1268156 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3ce, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ef, 10'h18c, 14'h00cf};
#1268160 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1268560 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3d5, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h154, 10'h18c, 14'h00c4};
#1268564 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1268964 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3db, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1b9, 10'h18c, 14'h00c9};
#1268968 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1269368 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3e1, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h21e, 10'h18c, 14'h00ce};
#1269372 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1269772 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3e8, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h283, 10'h18c, 14'h00c3};
#1269776 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1270176 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3ee, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2e8, 10'h18c, 14'h00c8};
#1270180 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1270580 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3c2, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02d, 10'h18d, 14'h00dd};
#1270584 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1270984 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3c9, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h092, 10'h18d, 14'h00d2};
#1270988 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1271388 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3cf, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0f7, 10'h18d, 14'h00d7};
#1271392 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1271792 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3d5, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h15c, 10'h18d, 14'h00dc};
#1271796 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1272196 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3dc, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1c1, 10'h18d, 14'h00d1};
#1272200 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1272600 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3e2, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h226, 10'h18d, 14'h00d6};
#1272604 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1273004 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3e8, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h28b, 10'h18d, 14'h00db};
#1273008 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1273408 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3ef, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2f0, 10'h18d, 14'h00d0};
#1273412 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1273812 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3c3, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h035, 10'h18e, 14'h00e5};
#1273816 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1274216 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3c9, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h09a, 10'h18e, 14'h00ea};
#1274220 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1274620 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3cf, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ff, 10'h18e, 14'h00ef};
#1274624 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1275024 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3d6, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h164, 10'h18e, 14'h00e4};
#1275028 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1275428 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3dc, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1c9, 10'h18e, 14'h00e9};
#1275432 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1275832 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3e2, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h22e, 10'h18e, 14'h00ee};
#1275836 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1276236 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3e9, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h293, 10'h18e, 14'h00e3};
#1276240 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1276640 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h3ef, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2f8, 10'h18e, 14'h00e8};
#1276644 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1357844 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h420, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h105, 10'h1a8, 14'h0085};
#1357848 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1358248 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h426, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h16a, 10'h1a8, 14'h008a};
#1358252 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1358652 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h42c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1cf, 10'h1a8, 14'h008f};
#1358656 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1359056 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h433, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h234, 10'h1a8, 14'h0084};
#1359060 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1359460 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h439, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h299, 10'h1a8, 14'h0089};
#1359464 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1359864 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h43f, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2fe, 10'h1a8, 14'h008e};
#1359868 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1360268 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h414, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h043, 10'h1a9, 14'h0093};
#1360272 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1360672 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h41a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0a8, 10'h1a9, 14'h0098};
#1360676 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1361076 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h420, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h10d, 10'h1a9, 14'h009d};
#1361080 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1361480 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h427, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h172, 10'h1a9, 14'h0092};
#1361484 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1361884 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h42d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1d7, 10'h1a9, 14'h0097};
#1361888 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1362288 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h433, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h23c, 10'h1a9, 14'h009c};
#1362292 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1362692 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h43a, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2a1, 10'h1a9, 14'h0091};
#1362696 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1363096 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h440, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h306, 10'h1a9, 14'h0096};
#1363100 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1363500 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h414, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h04b, 10'h1aa, 14'h00ab};
#1363504 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1363904 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h41b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0b0, 10'h1aa, 14'h00a0};
#1363908 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1364308 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h421, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h115, 10'h1aa, 14'h00a5};
#1364312 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1364712 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h427, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h17a, 10'h1aa, 14'h00aa};
#1364716 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1365116 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h42d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1df, 10'h1aa, 14'h00af};
#1365120 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1365520 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h434, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h244, 10'h1aa, 14'h00a4};
#1365524 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1365924 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h43a, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2a9, 10'h1aa, 14'h00a9};
#1365928 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1366328 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h440, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h30e, 10'h1aa, 14'h00ae};
#1366332 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1366732 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h415, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h053, 10'h1ab, 14'h00b3};
#1366736 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1367136 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h41b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0b8, 10'h1ab, 14'h00b8};
#1367140 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1367540 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h421, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h11d, 10'h1ab, 14'h00bd};
#1367544 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1367944 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h428, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h182, 10'h1ab, 14'h00b2};
#1367948 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1368348 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h42e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1e7, 10'h1ab, 14'h00b7};
#1368352 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1368752 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h434, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h24c, 10'h1ab, 14'h00bc};
#1368756 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1369156 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h43b, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2b1, 10'h1ab, 14'h00b1};
#1369160 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1369560 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h441, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h316, 10'h1ab, 14'h00b6};
#1369564 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1369964 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h415, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h05b, 10'h1ac, 14'h00cb};
#1369968 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1370368 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h41c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c0, 10'h1ac, 14'h00c0};
#1370372 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1370772 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h422, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h125, 10'h1ac, 14'h00c5};
#1370776 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1371176 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h428, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h18a, 10'h1ac, 14'h00ca};
#1371180 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1371580 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h42e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1ef, 10'h1ac, 14'h00cf};
#1371584 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1371984 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h435, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h254, 10'h1ac, 14'h00c4};
#1371988 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1372388 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h43b, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2b9, 10'h1ac, 14'h00c9};
#1372392 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1372792 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h441, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h31e, 10'h1ac, 14'h00ce};
#1372796 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1373196 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h416, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h063, 10'h1ad, 14'h00d3};
#1373200 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1373600 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h41c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c8, 10'h1ad, 14'h00d8};
#1373604 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1374004 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h422, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h12d, 10'h1ad, 14'h00dd};
#1374008 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1374408 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h429, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h192, 10'h1ad, 14'h00d2};
#1374412 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1374812 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h42f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1f7, 10'h1ad, 14'h00d7};
#1374816 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1375216 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h435, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h25c, 10'h1ad, 14'h00dc};
#1375220 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1375620 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h43c, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2c1, 10'h1ad, 14'h00d1};
#1375624 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1376024 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h410, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h006, 10'h1ae, 14'h00e6};
#1376028 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1376428 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h416, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h06b, 10'h1ae, 14'h00eb};
#1376432 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1376832 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h41d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d0, 10'h1ae, 14'h00e0};
#1376836 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1377236 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h423, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h135, 10'h1ae, 14'h00e5};
#1377240 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1377640 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h429, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h19a, 10'h1ae, 14'h00ea};
#1377644 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1458844 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h48c, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2c7, 10'h1c7, 14'h0077};
#1458848 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1459248 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h460, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00c, 10'h1c8, 14'h008c};
#1459252 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1459652 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h467, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h071, 10'h1c8, 14'h0081};
#1459656 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1460056 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h46d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d6, 10'h1c8, 14'h0086};
#1460060 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1460460 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h473, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h13b, 10'h1c8, 14'h008b};
#1460464 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1460864 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h47a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1a0, 10'h1c8, 14'h0080};
#1460868 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1461268 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h480, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h205, 10'h1c8, 14'h0085};
#1461272 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1461672 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h486, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h26a, 10'h1c8, 14'h008a};
#1461676 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1462076 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h48c, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2cf, 10'h1c8, 14'h008f};
#1462080 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1462480 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h461, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h014, 10'h1c9, 14'h0094};
#1462484 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1462884 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h467, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h079, 10'h1c9, 14'h0099};
#1462888 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1463288 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h46d, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0de, 10'h1c9, 14'h009e};
#1463292 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1463692 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h474, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h143, 10'h1c9, 14'h0093};
#1463696 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1464096 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h47a, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1a8, 10'h1c9, 14'h0098};
#1464100 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1464500 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h480, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h20d, 10'h1c9, 14'h009d};
#1464504 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1464904 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h487, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h272, 10'h1c9, 14'h0092};
#1464908 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1465308 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h48d, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2d7, 10'h1c9, 14'h0097};
#1465312 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1465712 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h461, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h01c, 10'h1ca, 14'h00ac};
#1465716 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1466116 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h468, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h081, 10'h1ca, 14'h00a1};
#1466120 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1466520 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h46e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e6, 10'h1ca, 14'h00a6};
#1466524 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1466924 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h474, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h14b, 10'h1ca, 14'h00ab};
#1466928 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1467328 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h47b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1b0, 10'h1ca, 14'h00a0};
#1467332 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1467732 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h481, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h215, 10'h1ca, 14'h00a5};
#1467736 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1468136 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h487, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h27a, 10'h1ca, 14'h00aa};
#1468140 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1468540 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h48d, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2df, 10'h1ca, 14'h00af};
#1468544 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1468944 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h462, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h024, 10'h1cb, 14'h00b4};
#1468948 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1469348 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h468, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h089, 10'h1cb, 14'h00b9};
#1469352 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1469752 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h46e, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ee, 10'h1cb, 14'h00be};
#1469756 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1470156 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h475, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h153, 10'h1cb, 14'h00b3};
#1470160 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1470560 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h47b, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1b8, 10'h1cb, 14'h00b8};
#1470564 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1470964 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h481, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h21d, 10'h1cb, 14'h00bd};
#1470968 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1471368 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h488, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h282, 10'h1cb, 14'h00b2};
#1471372 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1471772 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h48e, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2e7, 10'h1cb, 14'h00b7};
#1471776 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1472176 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h462, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02c, 10'h1cc, 14'h00cc};
#1472180 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1472580 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h469, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h091, 10'h1cc, 14'h00c1};
#1472584 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1472984 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h46f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0f6, 10'h1cc, 14'h00c6};
#1472988 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1473388 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h475, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h15b, 10'h1cc, 14'h00cb};
#1473392 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1473792 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h47c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1c0, 10'h1cc, 14'h00c0};
#1473796 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1474196 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h482, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h225, 10'h1cc, 14'h00c5};
#1474200 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1474600 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h488, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h28a, 10'h1cc, 14'h00ca};
#1474604 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1475004 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h48e, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2ef, 10'h1cc, 14'h00cf};
#1475008 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1475408 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h463, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h034, 10'h1cd, 14'h00d4};
#1475412 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1475812 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h469, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h099, 10'h1cd, 14'h00d9};
#1475816 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1476216 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h46f, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0fe, 10'h1cd, 14'h00de};
#1476220 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1476620 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h476, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h163, 10'h1cd, 14'h00d3};
#1476624 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1477024 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h47c, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h1c8, 10'h1cd, 14'h00d8};
#1477028 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1477428 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h482, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h22d, 10'h1cd, 14'h00dd};
#1477432 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1477832 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h489, 6'h00, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h292, 10'h1cd, 14'h00d2};
#1477836 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1478236 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h48f, 6'h00, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2f7, 10'h1cd, 14'h00d7};
#1478240 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1478640 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h463, 6'h00, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h03c, 10'h1ce, 14'h00ec};
#1478644 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1559844 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4c6, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h169, 10'h1e7, 14'hxx79};
#1559848 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1560248 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4cc, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h1ce, 10'h1e7, 14'hxx7e};
#1560252 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1560652 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4d3, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h233, 10'h1e7, 14'hxx73};
#1560656 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1561056 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4d9, 6'hxx, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h298, 10'h1e7, 14'hxx78};
#1561060 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1561460 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4df, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2fd, 10'h1e7, 14'hxx7d};
#1561464 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1561864 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4b4, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h042, 10'h1e8, 14'hxx82};
#1561868 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1562268 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4ba, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h0a7, 10'h1e8, 14'hxx87};
#1562272 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1562672 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4c0, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h10c, 10'h1e8, 14'hxx8c};
#1562676 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1563076 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4c7, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h171, 10'h1e8, 14'hxx81};
#1563080 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1563480 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4cd, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h1d6, 10'h1e8, 14'hxx86};
#1563484 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1563884 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4d3, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h23b, 10'h1e8, 14'hxx8b};
#1563888 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1564288 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4da, 6'hxx, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2a0, 10'h1e8, 14'hxx80};
#1564292 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1564692 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4e0, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h305, 10'h1e8, 14'hxx85};
#1564696 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1565096 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4b4, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h04a, 10'h1e9, 14'hxx9a};
#1565100 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1565500 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4ba, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h0af, 10'h1e9, 14'hxx9f};
#1565504 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1565904 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4c1, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h114, 10'h1e9, 14'hxx94};
#1565908 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1566308 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4c7, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h179, 10'h1e9, 14'hxx99};
#1566312 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1566712 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4cd, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h1de, 10'h1e9, 14'hxx9e};
#1566716 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1567116 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4d4, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h243, 10'h1e9, 14'hxx93};
#1567120 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1567520 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4da, 6'hxx, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2a8, 10'h1e9, 14'hxx98};
#1567524 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1567924 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4e0, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h30d, 10'h1e9, 14'hxx9d};
#1567928 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1568328 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4b5, 6'hxx, 1'b1, 1'b0, 4'h0, 4'h0, 4'h0, 10'h052, 10'h1ea, 14'hxxa2};
#1568332 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1568732 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4bb, 6'hxx, 1'b1, 1'b0, 4'h0, 4'h0, 4'h0, 10'h0b7, 10'h1ea, 14'hxxa7};
#1568736 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1569136 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4c1, 6'hxx, 1'b1, 1'b0, 4'h0, 4'h0, 4'h0, 10'h11c, 10'h1ea, 14'hxxac};
#1569140 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1569540 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4c8, 6'hxx, 1'b1, 1'b0, 4'h0, 4'h0, 4'h0, 10'h181, 10'h1ea, 14'hxxa1};
#1569544 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1569944 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4ce, 6'hxx, 1'b1, 1'b0, 4'h0, 4'h0, 4'h0, 10'h1e6, 10'h1ea, 14'hxxa6};
#1569948 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1570348 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4d4, 6'hxx, 1'b1, 1'b0, 4'h0, 4'h0, 4'h0, 10'h24b, 10'h1ea, 14'hxxab};
#1570352 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1570752 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4db, 6'hxx, 1'b0, 1'b0, 4'h0, 4'h0, 4'h0, 10'h2b0, 10'h1ea, 14'hxxa0};
#1570756 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1571156 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4e1, 6'hxx, 1'b1, 1'b0, 4'h0, 4'h0, 4'h0, 10'h315, 10'h1ea, 14'hxxa5};
#1571160 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1571560 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4b5, 6'hxx, 1'b1, 1'b0, 4'h0, 4'h0, 4'h0, 10'h05a, 10'h1eb, 14'hxxba};
#1571564 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1571964 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4bb, 6'hxx, 1'b1, 1'b0, 4'h0, 4'h0, 4'h0, 10'h0bf, 10'h1eb, 14'hxxbf};
#1571968 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1572368 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4c2, 6'hxx, 1'b1, 1'b0, 4'h0, 4'h0, 4'h0, 10'h124, 10'h1eb, 14'hxxb4};
#1572372 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1572772 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4c8, 6'hxx, 1'b1, 1'b0, 4'h0, 4'h0, 4'h0, 10'h189, 10'h1eb, 14'hxxb9};
#1572776 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1573176 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4ce, 6'hxx, 1'b1, 1'b0, 4'h0, 4'h0, 4'h0, 10'h1ee, 10'h1eb, 14'hxxbe};
#1573180 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1573580 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4d5, 6'hxx, 1'b1, 1'b0, 4'h0, 4'h0, 4'h0, 10'h253, 10'h1eb, 14'hxxb3};
#1573584 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1573984 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4db, 6'hxx, 1'b0, 1'b0, 4'h0, 4'h0, 4'h0, 10'h2b8, 10'h1eb, 14'hxxb8};
#1573988 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1574388 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4e1, 6'hxx, 1'b1, 1'b0, 4'h0, 4'h0, 4'h0, 10'h31d, 10'h1eb, 14'hxxbd};
#1574392 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1574792 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4b6, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h062, 10'h1ec, 14'hxxc2};
#1574796 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1575196 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4bc, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h0c7, 10'h1ec, 14'hxxc7};
#1575200 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1575600 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4c2, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h12c, 10'h1ec, 14'hxxcc};
#1575604 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1576004 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4c9, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h191, 10'h1ec, 14'hxxc1};
#1576008 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1576408 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4cf, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h1f6, 10'h1ec, 14'hxxc6};
#1576412 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1576812 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4d5, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h25b, 10'h1ec, 14'hxxcb};
#1576816 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1577216 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4dc, 6'hxx, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2c0, 10'h1ec, 14'hxxc0};
#1577220 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1577620 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4b0, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h005, 10'h1ed, 14'hxxd5};
#1577624 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1578024 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4b6, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h06a, 10'h1ed, 14'hxxda};
#1578028 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1578428 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4bc, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h0cf, 10'h1ed, 14'hxxdf};
#1578432 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1578832 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4c3, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h134, 10'h1ed, 14'hxxd4};
#1578836 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1579236 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4c9, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h199, 10'h1ed, 14'hxxd9};
#1579240 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1579640 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h4cf, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h1fe, 10'h1ed, 14'hxxde};
#1579644 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1660844 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h500, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h00b, 10'h207, 14'hxx7b};
#1660848 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1661248 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h507, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h070, 10'h207, 14'hxx70};
#1661252 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1661652 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h50d, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h0d5, 10'h207, 14'hxx75};
#1661656 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1662056 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h513, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h13a, 10'h207, 14'hxx7a};
#1662060 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1662460 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h519, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h19f, 10'h207, 14'hxx7f};
#1662464 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1662864 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h520, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h204, 10'h207, 14'hxx74};
#1662868 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1663268 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h526, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h269, 10'h207, 14'hxx79};
#1663272 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1663672 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h52c, 6'hxx, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2ce, 10'h207, 14'hxx7e};
#1663676 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1664076 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h501, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h013, 10'h208, 14'hxx83};
#1664080 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1664480 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h507, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h078, 10'h208, 14'hxx88};
#1664484 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1664884 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h50d, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h0dd, 10'h208, 14'hxx8d};
#1664888 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1665288 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h514, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h142, 10'h208, 14'hxx82};
#1665292 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1665692 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h51a, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h1a7, 10'h208, 14'hxx87};
#1665696 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1666096 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h520, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h20c, 10'h208, 14'hxx8c};
#1666100 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1666500 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h527, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h271, 10'h208, 14'hxx81};
#1666504 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1666904 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h52d, 6'hxx, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2d6, 10'h208, 14'hxx86};
#1666908 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1667308 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h501, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h01b, 10'h209, 14'hxx9b};
#1667312 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1667712 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h508, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h080, 10'h209, 14'hxx90};
#1667716 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1668116 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h50e, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h0e5, 10'h209, 14'hxx95};
#1668120 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1668520 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h514, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h14a, 10'h209, 14'hxx9a};
#1668524 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1668924 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h51a, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h1af, 10'h209, 14'hxx9f};
#1668928 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1669328 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h521, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h214, 10'h209, 14'hxx94};
#1669332 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1669732 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h527, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h279, 10'h209, 14'hxx99};
#1669736 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1670136 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h52d, 6'hxx, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2de, 10'h209, 14'hxx9e};
#1670140 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1670540 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h502, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h023, 10'h20a, 14'hxxa3};
#1670544 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1670944 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h508, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h088, 10'h20a, 14'hxxa8};
#1670948 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1671348 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h50e, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h0ed, 10'h20a, 14'hxxad};
#1671352 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1671752 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h515, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h152, 10'h20a, 14'hxxa2};
#1671756 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1672156 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h51b, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h1b7, 10'h20a, 14'hxxa7};
#1672160 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1672560 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h521, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h21c, 10'h20a, 14'hxxac};
#1672564 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1672964 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h528, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h281, 10'h20a, 14'hxxa1};
#1672968 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1673368 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h52e, 6'hxx, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2e6, 10'h20a, 14'hxxa6};
#1673372 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1673772 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h502, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h02b, 10'h20b, 14'hxxbb};
#1673776 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1674176 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h509, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h090, 10'h20b, 14'hxxb0};
#1674180 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1674580 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h50f, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h0f5, 10'h20b, 14'hxxb5};
#1674584 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1674984 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h515, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h15a, 10'h20b, 14'hxxba};
#1674988 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1675388 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h51b, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h1bf, 10'h20b, 14'hxxbf};
#1675392 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1675792 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h522, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h224, 10'h20b, 14'hxxb4};
#1675796 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1676196 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h528, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h289, 10'h20b, 14'hxxb9};
#1676200 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1676600 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h52e, 6'hxx, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2ee, 10'h20b, 14'hxxbe};
#1676604 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1677004 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h503, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h033, 10'h20c, 14'hxxc3};
#1677008 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1677408 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h509, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h098, 10'h20c, 14'hxxc8};
#1677412 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1677812 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h50f, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h0fd, 10'h20c, 14'hxxcd};
#1677816 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1678216 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h516, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h162, 10'h20c, 14'hxxc2};
#1678220 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1678620 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h51c, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h1c7, 10'h20c, 14'hxxc7};
#1678624 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1679024 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h522, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h22c, 10'h20c, 14'hxxcc};
#1679028 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1679428 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h529, 6'hxx, 1'b0, 1'b1, 4'h0, 4'h0, 4'h0, 10'h291, 10'h20c, 14'hxxc1};
#1679432 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};
#1679832 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr} <= {11'h52f, 6'hxx, 1'b1, 1'b1, 4'h0, 4'h0, 4'h0, 10'h2f6, 10'h20c, 14'hxxc6};
#1679836 {smem_addr, charcode, hsync, vsync, red, green, blue, x, y, bmem_addr}  <= {65{1'b x}};


join
end

endmodule